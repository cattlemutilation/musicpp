----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date:    14:24:35 10/08/2019 
-- Design Name: 
-- Module Name:    rom - Behavioral 
-- Project Name: 
-- Target Devices: 
-- Tool versions: 
-- Description: 
--
-- Dependencies: 
--
-- Revision: 
-- Revision 0.01 - File Created
-- Additional Comments: 
--
----------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--use IEEE.NUMERIC_STD.ALL;

-- Uncomment the following library declaration if instantiating
-- any Xilinx primitives in this code.
--library UNISIM;
--use UNISIM.VComponents.all;

--named rom but is actually ram
entity ram is
    Port ( clk : in  STD_LOGIC;
           rst : in  STD_LOGIC;
			  wr_en : in STD_LOGIC;
           addr : in  STD_LOGIC_VECTOR (10 downto 0);
			  data_in : in STD_LOGIC_VECTOR(7 downto 0);
           data_out : out  STD_LOGIC_VECTOR (7 downto 0));
end rom;

architecture Behavioral of ram is

type ram_type is array (2047 downto 0) of std_logic_vector(7 downto 0);
signal ram : ram_type;

begin

	ram_process: process(clk, addr) is
	variable var_ram : ram_type;
	variable var_addr : integer;
	
	begin
		if (rst = '1') then
		
		var_ram(0) := "00000001";
		var_ram(1) := "00000001";
		var_ram(2) := "00111100";	-- start
		var_ram(3) := "00000001";	-- semiquaver
		var_ram(4) := "01110001";	-- e5
		var_ram(5) := "00000001";	-- semiq
		var_ram(6) := "01110000";	-- d5#
		var_ram(7) := "00000001"; 
		var_ram(8) := "01110001"; -- e5
		var_ram(9) := "00000001"; 
		var_ram(10) := "01110000"; -- d5#
		var_ram(11) := "00000001";
		var_ram(12) := "01110001"; -- e5
		var_ram(13) := "00000001";
		var_ram(14) := "01101100"; -- b4
		var_ram(15) := "00000001";
		var_ram(16) := "01101111"; -- d5
		var_ram(17) := "00000001";	
		var_ram(18) := "01101101"; -- c5
		var_ram(19) := "00000010";-- quaver
		var_ram(20) := "01101010"; -- a4
		var_ram(21) := "00000001";
		var_ram(22) := "00000000"; -- resti  guess
		var_ram(23) := "00000001"; 
		var_ram(24) := "01100001";
		var_ram(25) := "00000001";
		var_ram(26) := "01100101";
		var_ram(27) := "00000001";
		var_ram(28) := "01101010";
		var_ram(29) := "00000010";
		var_ram(30) := "01101100"; -- b4
		var_ram(31) := "00000001";
		var_ram(32) := "00000000"; -- rest
		var_ram(33) := "00000001";
		var_ram(34) := "01100101"; -- e
		var_ram(35) := "00000001";
		var_ram(36) := "01101001"; -- g#
		var_ram(37) := "00000001";
		var_ram(38) := "01101100"; -- b
		var_ram(39) := "00000010";
		var_ram(40) := "01101101"; -- c
		var_ram(41) := "00000001"; 
		var_ram(42) := "00000000";
		var_ram(43) := "01000000";
		var_ram(44) := "00000000";
		var_ram(45) := "00000000";
		var_ram(46) := "00000000";
		var_ram(47) := "00000000";
		var_ram(48) := "00000000";
		var_ram(49) := "00000000";
		var_ram(50) := "00000000";
		var_ram(51) := "00000000";
		var_ram(52) := "00000000";
		var_ram(53) := "00000000";
		var_ram(54) := "00000000";
		var_ram(55) := "00000000";
		var_ram(56) := "00000000";
		var_ram(57) := "00000000";
		var_ram(58) := "00000000";
		var_ram(59) := "00000000";
		var_ram(60) := "00000000";
		var_ram(61) := "00000000";
		var_ram(62) := "00000000";
		var_ram(63) := "00000000";
		var_ram(64) := "00000000";
		var_ram(65) := "00000000";
		var_ram(66) := "00000000";
		var_ram(67) := "00000000";
		var_ram(68) := "00000000";
		var_ram(69) := "00000000";
		var_ram(70) := "00000000";
		var_ram(71) := "00000000";
		var_ram(72) := "00000000";
		var_ram(73) := "00000000";
		var_ram(74) := "00000000";
		var_ram(75) := "00000000";
		var_ram(76) := "00000000";
		var_ram(77) := "00000000";
		var_ram(78) := "00000000";
		var_ram(79) := "00000000";
		var_ram(80) := "00000000";
		var_ram(81) := "00000000";
		var_ram(82) := "00000000";
		var_ram(83) := "00000000";
		var_ram(84) := "00000000";
		var_ram(85) := "00000000";
		var_ram(86) := "00000000";
		var_ram(87) := "00000000";
		var_ram(88) := "00000000";
		var_ram(89) := "00000000";
		var_ram(90) := "00000000";
		var_ram(91) := "00000000";
		var_ram(92) := "00000000";
		var_ram(93) := "00000000";
		var_ram(94) := "00000000";
		var_ram(95) := "00000000";
		var_ram(96) := "00000000";
		var_ram(97) := "00000000";
		var_ram(98) := "00000000";
		var_ram(99) := "00000000";
		var_ram(100) := "00000000";
		var_ram(101) := "00000000";
		var_ram(102) := "00000000";
		var_ram(103) := "00000000";
		var_ram(104) := "00000000";
		var_ram(105) := "00000000";
		var_ram(106) := "00000000";
		var_ram(107) := "00000000";
		var_ram(108) := "00000000";
		var_ram(109) := "00000000";
		var_ram(110) := "00000000";
		var_ram(111) := "00000000";
		var_ram(112) := "00000000";
		var_ram(113) := "00000000";
		var_ram(114) := "00000000";
		var_ram(115) := "00000000";
		var_ram(116) := "00000000";
		var_ram(117) := "00000000";
		var_ram(118) := "00000000";
		var_ram(119) := "00000000";
		var_ram(120) := "00000000";
		var_ram(121) := "00000000";
		var_ram(122) := "00000000";
		var_ram(123) := "00000000";
		var_ram(124) := "00000000";
		var_ram(125) := "00000000";
		var_ram(126) := "00000000";
		var_ram(127) := "00000000";
		var_ram(128) := "00000000";
		var_ram(129) := "00000000";
		var_ram(130) := "00000000";
		var_ram(131) := "00000000";
		var_ram(132) := "00000000";
		var_ram(133) := "00000000";
		var_ram(134) := "00000000";
		var_ram(135) := "00000000";
		var_ram(136) := "00000000";
		var_ram(137) := "00000000";
		var_ram(138) := "00000000";
		var_ram(139) := "00000000";
		var_ram(140) := "00000000";
		var_ram(141) := "00000000";
		var_ram(142) := "00000000";
		var_ram(143) := "00000000";
		var_ram(144) := "00000000";
		var_ram(145) := "00000000";
		var_ram(146) := "00000000";
		var_ram(147) := "00000000";
		var_ram(148) := "00000000";
		var_ram(149) := "00000000";
		var_ram(150) := "00000000";
		var_ram(151) := "00000000";
		var_ram(152) := "00000000";
		var_ram(153) := "00000000";
		var_ram(154) := "00000000";
		var_ram(155) := "00000000";
		var_ram(156) := "00000000";
		var_ram(157) := "00000000";
		var_ram(158) := "00000000";
		var_ram(159) := "00000000";
		var_ram(160) := "00000000";
		var_ram(161) := "00000000";
		var_ram(162) := "00000000";
		var_ram(163) := "00000000";
		var_ram(164) := "00000000";
		var_ram(165) := "00000000";
		var_ram(166) := "00000000";
		var_ram(167) := "00000000";
		var_ram(168) := "00000000";
		var_ram(169) := "00000000";
		var_ram(170) := "00000000";
		var_ram(171) := "00000000";
		var_ram(172) := "00000000";
		var_ram(173) := "00000000";
		var_ram(174) := "00000000";
		var_ram(175) := "00000000";
		var_ram(176) := "00000000";
		var_ram(177) := "00000000";
		var_ram(178) := "00000000";
		var_ram(179) := "00000000";
		var_ram(180) := "00000000";
		var_ram(181) := "00000000";
		var_ram(182) := "00000000";
		var_ram(183) := "00000000";
		var_ram(184) := "00000000";
		var_ram(185) := "00000000";
		var_ram(186) := "00000000";
		var_ram(187) := "00000000";
		var_ram(188) := "00000000";
		var_ram(189) := "00000000";
		var_ram(190) := "00000000";
		var_ram(191) := "00000000";
		var_ram(192) := "00000000";
		var_ram(193) := "00000000";
		var_ram(194) := "00000000";
		var_ram(195) := "00000000";
		var_ram(196) := "00000000";
		var_ram(197) := "00000000";
		var_ram(198) := "00000000";
		var_ram(199) := "00000000";
		var_ram(200) := "00000000";
		var_ram(201) := "00000000";
		var_ram(202) := "00000000";
		var_ram(203) := "00000000";
		var_ram(204) := "00000000";
		var_ram(205) := "00000000";
		var_ram(206) := "00000000";
		var_ram(207) := "00000000";
		var_ram(208) := "00000000";
		var_ram(209) := "00000000";
		var_ram(210) := "00000000";
		var_ram(211) := "00000000";
		var_ram(212) := "00000000";
		var_ram(213) := "00000000";
		var_ram(214) := "00000000";
		var_ram(215) := "00000000";
		var_ram(216) := "00000000";
		var_ram(217) := "00000000";
		var_ram(218) := "00000000";
		var_ram(219) := "00000000";
		var_ram(220) := "00000000";
		var_ram(221) := "00000000";
		var_ram(222) := "00000000";
		var_ram(223) := "00000000";
		var_ram(224) := "00000000";
		var_ram(225) := "00000000";
		var_ram(226) := "00000000";
		var_ram(227) := "00000000";
		var_ram(228) := "00000000";
		var_ram(229) := "00000000";
		var_ram(230) := "00000000";
		var_ram(231) := "00000000";
		var_ram(232) := "00000000";
		var_ram(233) := "00000000";
		var_ram(234) := "00000000";
		var_ram(235) := "00000000";
		var_ram(236) := "00000000";
		var_ram(237) := "00000000";
		var_ram(238) := "00000000";
		var_ram(239) := "00000000";
		var_ram(240) := "00000000";
		var_ram(241) := "00000000";
		var_ram(242) := "00000000";
		var_ram(243) := "00000000";
		var_ram(244) := "00000000";
		var_ram(245) := "00000000";
		var_ram(246) := "00000000";
		var_ram(247) := "00000000";
		var_ram(248) := "00000000";
		var_ram(249) := "00000000";
		var_ram(250) := "00000000";
		var_ram(251) := "00000000";
		var_ram(252) := "00000000";
		var_ram(253) := "00000000";
		var_ram(254) := "00000000";
		var_ram(255) := "00000000";
		var_ram(256) := "00000000";
		var_ram(257) := "00000000";
		var_ram(258) := "00000000";
		var_ram(259) := "00000000";
		var_ram(260) := "00000000";
		var_ram(261) := "00000000";
		var_ram(262) := "00000000";
		var_ram(263) := "00000000";
		var_ram(264) := "00000000";
		var_ram(265) := "00000000";
		var_ram(266) := "00000000";
		var_ram(267) := "00000000";
		var_ram(268) := "00000000";
		var_ram(269) := "00000000";
		var_ram(270) := "00000000";
		var_ram(271) := "00000000";
		var_ram(272) := "00000000";
		var_ram(273) := "00000000";
		var_ram(274) := "00000000";
		var_ram(275) := "00000000";
		var_ram(276) := "00000000";
		var_ram(277) := "00000000";
		var_ram(278) := "00000000";
		var_ram(279) := "00000000";
		var_ram(280) := "00000000";
		var_ram(281) := "00000000";
		var_ram(282) := "00000000";
		var_ram(283) := "00000000";
		var_ram(284) := "00000000";
		var_ram(285) := "00000000";
		var_ram(286) := "00000000";
		var_ram(287) := "00000000";
		var_ram(288) := "00000000";
		var_ram(289) := "00000000";
		var_ram(290) := "00000000";
		var_ram(291) := "00000000";
		var_ram(292) := "00000000";
		var_ram(293) := "00000000";
		var_ram(294) := "00000000";
		var_ram(295) := "00000000";
		var_ram(296) := "00000000";
		var_ram(297) := "00000000";
		var_ram(298) := "00000000";
		var_ram(299) := "00000000";
		var_ram(300) := "00000000";
		var_ram(301) := "00000000";
		var_ram(302) := "00000000";
		var_ram(303) := "00000000";
		var_ram(304) := "00000000";
		var_ram(305) := "00000000";
		var_ram(306) := "00000000";
		var_ram(307) := "00000000";
		var_ram(308) := "00000000";
		var_ram(309) := "00000000";
		var_ram(310) := "00000000";
		var_ram(311) := "00000000";
		var_ram(312) := "00000000";
		var_ram(313) := "00000000";
		var_ram(314) := "00000000";
		var_ram(315) := "00000000";
		var_ram(316) := "00000000";
		var_ram(317) := "00000000";
		var_ram(318) := "00000000";
		var_ram(319) := "00000000";
		var_ram(320) := "00000000";
		var_ram(321) := "00000000";
		var_ram(322) := "00000000";
		var_ram(323) := "00000000";
		var_ram(324) := "00000000";
		var_ram(325) := "00000000";
		var_ram(326) := "00000000";
		var_ram(327) := "00000000";
		var_ram(328) := "00000000";
		var_ram(329) := "00000000";
		var_ram(330) := "00000000";
		var_ram(331) := "00000000";
		var_ram(332) := "00000000";
		var_ram(333) := "00000000";
		var_ram(334) := "00000000";
		var_ram(335) := "00000000";
		var_ram(336) := "00000000";
		var_ram(337) := "00000000";
		var_ram(338) := "00000000";
		var_ram(339) := "00000000";
		var_ram(340) := "00000000";
		var_ram(341) := "00000000";
		var_ram(342) := "00000000";
		var_ram(343) := "00000000";
		var_ram(344) := "00000000";
		var_ram(345) := "00000000";
		var_ram(346) := "00000000";
		var_ram(347) := "00000000";
		var_ram(348) := "00000000";
		var_ram(349) := "00000000";
		var_ram(350) := "00000000";
		var_ram(351) := "00000000";
		var_ram(352) := "00000000";
		var_ram(353) := "00000000";
		var_ram(354) := "00000000";
		var_ram(355) := "00000000";
		var_ram(356) := "00000000";
		var_ram(357) := "00000000";
		var_ram(358) := "00000000";
		var_ram(359) := "00000000";
		var_ram(360) := "00000000";
		var_ram(361) := "00000000";
		var_ram(362) := "00000000";
		var_ram(363) := "00000000";
		var_ram(364) := "00000000";
		var_ram(365) := "00000000";
		var_ram(366) := "00000000";
		var_ram(367) := "00000000";
		var_ram(368) := "00000000";
		var_ram(369) := "00000000";
		var_ram(370) := "00000000";
		var_ram(371) := "00000000";
		var_ram(372) := "00000000";
		var_ram(373) := "00000000";
		var_ram(374) := "00000000";
		var_ram(375) := "00000000";
		var_ram(376) := "00000000";
		var_ram(377) := "00000000";
		var_ram(378) := "00000000";
		var_ram(379) := "00000000";
		var_ram(380) := "00000000";
		var_ram(381) := "00000000";
		var_ram(382) := "00000000";
		var_ram(383) := "00000000";
		var_ram(384) := "00000000";
		var_ram(385) := "00000000";
		var_ram(386) := "00000000";
		var_ram(387) := "00000000";
		var_ram(388) := "00000000";
		var_ram(389) := "00000000";
		var_ram(390) := "00000000";
		var_ram(391) := "00000000";
		var_ram(392) := "00000000";
		var_ram(393) := "00000000";
		var_ram(394) := "00000000";
		var_ram(395) := "00000000";
		var_ram(396) := "00000000";
		var_ram(397) := "00000000";
		var_ram(398) := "00000000";
		var_ram(399) := "00000000";
		var_ram(400) := "00000000";
		var_ram(401) := "00000000";
		var_ram(402) := "00000000";
		var_ram(403) := "00000000";
		var_ram(404) := "00000000";
		var_ram(405) := "00000000";
		var_ram(406) := "00000000";
		var_ram(407) := "00000000";
		var_ram(408) := "00000000";
		var_ram(409) := "00000000";
		var_ram(410) := "00000000";
		var_ram(411) := "00000000";
		var_ram(412) := "00000000";
		var_ram(413) := "00000000";
		var_ram(414) := "00000000";
		var_ram(415) := "00000000";
		var_ram(416) := "00000000";
		var_ram(417) := "00000000";
		var_ram(418) := "00000000";
		var_ram(419) := "00000000";
		var_ram(420) := "00000000";
		var_ram(421) := "00000000";
		var_ram(422) := "00000000";
		var_ram(423) := "00000000";
		var_ram(424) := "00000000";
		var_ram(425) := "00000000";
		var_ram(426) := "00000000";
		var_ram(427) := "00000000";
		var_ram(428) := "00000000";
		var_ram(429) := "00000000";
		var_ram(430) := "00000000";
		var_ram(431) := "00000000";
		var_ram(432) := "00000000";
		var_ram(433) := "00000000";
		var_ram(434) := "00000000";
		var_ram(435) := "00000000";
		var_ram(436) := "00000000";
		var_ram(437) := "00000000";
		var_ram(438) := "00000000";
		var_ram(439) := "00000000";
		var_ram(440) := "00000000";
		var_ram(441) := "00000000";
		var_ram(442) := "00000000";
		var_ram(443) := "00000000";
		var_ram(444) := "00000000";
		var_ram(445) := "00000000";
		var_ram(446) := "00000000";
		var_ram(447) := "00000000";
		var_ram(448) := "00000000";
		var_ram(449) := "00000000";
		var_ram(450) := "00000000";
		var_ram(451) := "00000000";
		var_ram(452) := "00000000";
		var_ram(453) := "00000000";
		var_ram(454) := "00000000";
		var_ram(455) := "00000000";
		var_ram(456) := "00000000";
		var_ram(457) := "00000000";
		var_ram(458) := "00000000";
		var_ram(459) := "00000000";
		var_ram(460) := "00000000";
		var_ram(461) := "00000000";
		var_ram(462) := "00000000";
		var_ram(463) := "00000000";
		var_ram(464) := "00000000";
		var_ram(465) := "00000000";
		var_ram(466) := "00000000";
		var_ram(467) := "00000000";
		var_ram(468) := "00000000";
		var_ram(469) := "00000000";
		var_ram(470) := "00000000";
		var_ram(471) := "00000000";
		var_ram(472) := "00000000";
		var_ram(473) := "00000000";
		var_ram(474) := "00000000";
		var_ram(475) := "00000000";
		var_ram(476) := "00000000";
		var_ram(477) := "00000000";
		var_ram(478) := "00000000";
		var_ram(479) := "00000000";
		var_ram(480) := "00000000";
		var_ram(481) := "00000000";
		var_ram(482) := "00000000";
		var_ram(483) := "00000000";
		var_ram(484) := "00000000";
		var_ram(485) := "00000000";
		var_ram(486) := "00000000";
		var_ram(487) := "00000000";
		var_ram(488) := "00000000";
		var_ram(489) := "00000000";
		var_ram(490) := "00000000";
		var_ram(491) := "00000000";
		var_ram(492) := "00000000";
		var_ram(493) := "00000000";
		var_ram(494) := "00000000";
		var_ram(495) := "00000000";
		var_ram(496) := "00000000";
		var_ram(497) := "00000000";
		var_ram(498) := "00000000";
		var_ram(499) := "00000000";
		var_ram(500) := "00000000";
		var_ram(501) := "00000000";
		var_ram(502) := "00000000";
		var_ram(503) := "00000000";
		var_ram(504) := "00000000";
		var_ram(505) := "00000000";
		var_ram(506) := "00000000";
		var_ram(507) := "00000000";
		var_ram(508) := "00000000";
		var_ram(509) := "00000000";
		var_ram(510) := "00000000";
		var_ram(511) := "00000000";
		var_ram(512) := "00000000";
		var_ram(513) := "00000000";
		var_ram(514) := "00000000";
		var_ram(515) := "00000000";
		var_ram(516) := "00000000";
		var_ram(517) := "00000000";
		var_ram(518) := "00000000";
		var_ram(519) := "00000000";
		var_ram(520) := "00000000";
		var_ram(521) := "00000000";
		var_ram(522) := "00000000";
		var_ram(523) := "00000000";
		var_ram(524) := "00000000";
		var_ram(525) := "00000000";
		var_ram(526) := "00000000";
		var_ram(527) := "00000000";
		var_ram(528) := "00000000";
		var_ram(529) := "00000000";
		var_ram(530) := "00000000";
		var_ram(531) := "00000000";
		var_ram(532) := "00000000";
		var_ram(533) := "00000000";
		var_ram(534) := "00000000";
		var_ram(535) := "00000000";
		var_ram(536) := "00000000";
		var_ram(537) := "00000000";
		var_ram(538) := "00000000";
		var_ram(539) := "00000000";
		var_ram(540) := "00000000";
		var_ram(541) := "00000000";
		var_ram(542) := "00000000";
		var_ram(543) := "00000000";
		var_ram(544) := "00000000";
		var_ram(545) := "00000000";
		var_ram(546) := "00000000";
		var_ram(547) := "00000000";
		var_ram(548) := "00000000";
		var_ram(549) := "00000000";
		var_ram(550) := "00000000";
		var_ram(551) := "00000000";
		var_ram(552) := "00000000";
		var_ram(553) := "00000000";
		var_ram(554) := "00000000";
		var_ram(555) := "00000000";
		var_ram(556) := "00000000";
		var_ram(557) := "00000000";
		var_ram(558) := "00000000";
		var_ram(559) := "00000000";
		var_ram(560) := "00000000";
		var_ram(561) := "00000000";
		var_ram(562) := "00000000";
		var_ram(563) := "00000000";
		var_ram(564) := "00000000";
		var_ram(565) := "00000000";
		var_ram(566) := "00000000";
		var_ram(567) := "00000000";
		var_ram(568) := "00000000";
		var_ram(569) := "00000000";
		var_ram(570) := "00000000";
		var_ram(571) := "00000000";
		var_ram(572) := "00000000";
		var_ram(573) := "00000000";
		var_ram(574) := "00000000";
		var_ram(575) := "00000000";
		var_ram(576) := "00000000";
		var_ram(577) := "00000000";
		var_ram(578) := "00000000";
		var_ram(579) := "00000000";
		var_ram(580) := "00000000";
		var_ram(581) := "00000000";
		var_ram(582) := "00000000";
		var_ram(583) := "00000000";
		var_ram(584) := "00000000";
		var_ram(585) := "00000000";
		var_ram(586) := "00000000";
		var_ram(587) := "00000000";
		var_ram(588) := "00000000";
		var_ram(589) := "00000000";
		var_ram(590) := "00000000";
		var_ram(591) := "00000000";
		var_ram(592) := "00000000";
		var_ram(593) := "00000000";
		var_ram(594) := "00000000";
		var_ram(595) := "00000000";
		var_ram(596) := "00000000";
		var_ram(597) := "00000000";
		var_ram(598) := "00000000";
		var_ram(599) := "00000000";
		var_ram(600) := "00000000";
		var_ram(601) := "00000000";
		var_ram(602) := "00000000";
		var_ram(603) := "00000000";
		var_ram(604) := "00000000";
		var_ram(605) := "00000000";
		var_ram(606) := "00000000";
		var_ram(607) := "00000000";
		var_ram(608) := "00000000";
		var_ram(609) := "00000000";
		var_ram(610) := "00000000";
		var_ram(611) := "00000000";
		var_ram(612) := "00000000";
		var_ram(613) := "00000000";
		var_ram(614) := "00000000";
		var_ram(615) := "00000000";
		var_ram(616) := "00000000";
		var_ram(617) := "00000000";
		var_ram(618) := "00000000";
		var_ram(619) := "00000000";
		var_ram(620) := "00000000";
		var_ram(621) := "00000000";
		var_ram(622) := "00000000";
		var_ram(623) := "00000000";
		var_ram(624) := "00000000";
		var_ram(625) := "00000000";
		var_ram(626) := "00000000";
		var_ram(627) := "00000000";
		var_ram(628) := "00000000";
		var_ram(629) := "00000000";
		var_ram(630) := "00000000";
		var_ram(631) := "00000000";
		var_ram(632) := "00000000";
		var_ram(633) := "00000000";
		var_ram(634) := "00000000";
		var_ram(635) := "00000000";
		var_ram(636) := "00000000";
		var_ram(637) := "00000000";
		var_ram(638) := "00000000";
		var_ram(639) := "00000000";
		var_ram(640) := "00000000";
		var_ram(641) := "00000000";
		var_ram(642) := "00000000";
		var_ram(643) := "00000000";
		var_ram(644) := "00000000";
		var_ram(645) := "00000000";
		var_ram(646) := "00000000";
		var_ram(647) := "00000000";
		var_ram(648) := "00000000";
		var_ram(649) := "00000000";
		var_ram(650) := "00000000";
		var_ram(651) := "00000000";
		var_ram(652) := "00000000";
		var_ram(653) := "00000000";
		var_ram(654) := "00000000";
		var_ram(655) := "00000000";
		var_ram(656) := "00000000";
		var_ram(657) := "00000000";
		var_ram(658) := "00000000";
		var_ram(659) := "00000000";
		var_ram(660) := "00000000";
		var_ram(661) := "00000000";
		var_ram(662) := "00000000";
		var_ram(663) := "00000000";
		var_ram(664) := "00000000";
		var_ram(665) := "00000000";
		var_ram(666) := "00000000";
		var_ram(667) := "00000000";
		var_ram(668) := "00000000";
		var_ram(669) := "00000000";
		var_ram(670) := "00000000";
		var_ram(671) := "00000000";
		var_ram(672) := "00000000";
		var_ram(673) := "00000000";
		var_ram(674) := "00000000";
		var_ram(675) := "00000000";
		var_ram(676) := "00000000";
		var_ram(677) := "00000000";
		var_ram(678) := "00000000";
		var_ram(679) := "00000000";
		var_ram(680) := "00000000";
		var_ram(681) := "00000000";
		var_ram(682) := "00000000";
		var_ram(683) := "00000000";
		var_ram(684) := "00000000";
		var_ram(685) := "00000000";
		var_ram(686) := "00000000";
		var_ram(687) := "00000000";
		var_ram(688) := "00000000";
		var_ram(689) := "00000000";
		var_ram(690) := "00000000";
		var_ram(691) := "00000000";
		var_ram(692) := "00000000";
		var_ram(693) := "00000000";
		var_ram(694) := "00000000";
		var_ram(695) := "00000000";
		var_ram(696) := "00000000";
		var_ram(697) := "00000000";
		var_ram(698) := "00000000";
		var_ram(699) := "00000000";
		var_ram(700) := "00000000";
		var_ram(701) := "00000000";
		var_ram(702) := "00000000";
		var_ram(703) := "00000000";
		var_ram(704) := "00000000";
		var_ram(705) := "00000000";
		var_ram(706) := "00000000";
		var_ram(707) := "00000000";
		var_ram(708) := "00000000";
		var_ram(709) := "00000000";
		var_ram(710) := "00000000";
		var_ram(711) := "00000000";
		var_ram(712) := "00000000";
		var_ram(713) := "00000000";
		var_ram(714) := "00000000";
		var_ram(715) := "00000000";
		var_ram(716) := "00000000";
		var_ram(717) := "00000000";
		var_ram(718) := "00000000";
		var_ram(719) := "00000000";
		var_ram(720) := "00000000";
		var_ram(721) := "00000000";
		var_ram(722) := "00000000";
		var_ram(723) := "00000000";
		var_ram(724) := "00000000";
		var_ram(725) := "00000000";
		var_ram(726) := "00000000";
		var_ram(727) := "00000000";
		var_ram(728) := "00000000";
		var_ram(729) := "00000000";
		var_ram(730) := "00000000";
		var_ram(731) := "00000000";
		var_ram(732) := "00000000";
		var_ram(733) := "00000000";
		var_ram(734) := "00000000";
		var_ram(735) := "00000000";
		var_ram(736) := "00000000";
		var_ram(737) := "00000000";
		var_ram(738) := "00000000";
		var_ram(739) := "00000000";
		var_ram(740) := "00000000";
		var_ram(741) := "00000000";
		var_ram(742) := "00000000";
		var_ram(743) := "00000000";
		var_ram(744) := "00000000";
		var_ram(745) := "00000000";
		var_ram(746) := "00000000";
		var_ram(747) := "00000000";
		var_ram(748) := "00000000";
		var_ram(749) := "00000000";
		var_ram(750) := "00000000";
		var_ram(751) := "00000000";
		var_ram(752) := "00000000";
		var_ram(753) := "00000000";
		var_ram(754) := "00000000";
		var_ram(755) := "00000000";
		var_ram(756) := "00000000";
		var_ram(757) := "00000000";
		var_ram(758) := "00000000";
		var_ram(759) := "00000000";
		var_ram(760) := "00000000";
		var_ram(761) := "00000000";
		var_ram(762) := "00000000";
		var_ram(763) := "00000000";
		var_ram(764) := "00000000";
		var_ram(765) := "00000000";
		var_ram(766) := "00000000";
		var_ram(767) := "00000000";
		var_ram(768) := "00000000";
		var_ram(769) := "00000000";
		var_ram(770) := "00000000";
		var_ram(771) := "00000000";
		var_ram(772) := "00000000";
		var_ram(773) := "00000000";
		var_ram(774) := "00000000";
		var_ram(775) := "00000000";
		var_ram(776) := "00000000";
		var_ram(777) := "00000000";
		var_ram(778) := "00000000";
		var_ram(779) := "00000000";
		var_ram(780) := "00000000";
		var_ram(781) := "00000000";
		var_ram(782) := "00000000";
		var_ram(783) := "00000000";
		var_ram(784) := "00000000";
		var_ram(785) := "00000000";
		var_ram(786) := "00000000";
		var_ram(787) := "00000000";
		var_ram(788) := "00000000";
		var_ram(789) := "00000000";
		var_ram(790) := "00000000";
		var_ram(791) := "00000000";
		var_ram(792) := "00000000";
		var_ram(793) := "00000000";
		var_ram(794) := "00000000";
		var_ram(795) := "00000000";
		var_ram(796) := "00000000";
		var_ram(797) := "00000000";
		var_ram(798) := "00000000";
		var_ram(799) := "00000000";
		var_ram(800) := "00000000";
		var_ram(801) := "00000000";
		var_ram(802) := "00000000";
		var_ram(803) := "00000000";
		var_ram(804) := "00000000";
		var_ram(805) := "00000000";
		var_ram(806) := "00000000";
		var_ram(807) := "00000000";
		var_ram(808) := "00000000";
		var_ram(809) := "00000000";
		var_ram(810) := "00000000";
		var_ram(811) := "00000000";
		var_ram(812) := "00000000";
		var_ram(813) := "00000000";
		var_ram(814) := "00000000";
		var_ram(815) := "00000000";
		var_ram(816) := "00000000";
		var_ram(817) := "00000000";
		var_ram(818) := "00000000";
		var_ram(819) := "00000000";
		var_ram(820) := "00000000";
		var_ram(821) := "00000000";
		var_ram(822) := "00000000";
		var_ram(823) := "00000000";
		var_ram(824) := "00000000";
		var_ram(825) := "00000000";
		var_ram(826) := "00000000";
		var_ram(827) := "00000000";
		var_ram(828) := "00000000";
		var_ram(829) := "00000000";
		var_ram(830) := "00000000";
		var_ram(831) := "00000000";
		var_ram(832) := "00000000";
		var_ram(833) := "00000000";
		var_ram(834) := "00000000";
		var_ram(835) := "00000000";
		var_ram(836) := "00000000";
		var_ram(837) := "00000000";
		var_ram(838) := "00000000";
		var_ram(839) := "00000000";
		var_ram(840) := "00000000";
		var_ram(841) := "00000000";
		var_ram(842) := "00000000";
		var_ram(843) := "00000000";
		var_ram(844) := "00000000";
		var_ram(845) := "00000000";
		var_ram(846) := "00000000";
		var_ram(847) := "00000000";
		var_ram(848) := "00000000";
		var_ram(849) := "00000000";
		var_ram(850) := "00000000";
		var_ram(851) := "00000000";
		var_ram(852) := "00000000";
		var_ram(853) := "00000000";
		var_ram(854) := "00000000";
		var_ram(855) := "00000000";
		var_ram(856) := "00000000";
		var_ram(857) := "00000000";
		var_ram(858) := "00000000";
		var_ram(859) := "00000000";
		var_ram(860) := "00000000";
		var_ram(861) := "00000000";
		var_ram(862) := "00000000";
		var_ram(863) := "00000000";
		var_ram(864) := "00000000";
		var_ram(865) := "00000000";
		var_ram(866) := "00000000";
		var_ram(867) := "00000000";
		var_ram(868) := "00000000";
		var_ram(869) := "00000000";
		var_ram(870) := "00000000";
		var_ram(871) := "00000000";
		var_ram(872) := "00000000";
		var_ram(873) := "00000000";
		var_ram(874) := "00000000";
		var_ram(875) := "00000000";
		var_ram(876) := "00000000";
		var_ram(877) := "00000000";
		var_ram(878) := "00000000";
		var_ram(879) := "00000000";
		var_ram(880) := "00000000";
		var_ram(881) := "00000000";
		var_ram(882) := "00000000";
		var_ram(883) := "00000000";
		var_ram(884) := "00000000";
		var_ram(885) := "00000000";
		var_ram(886) := "00000000";
		var_ram(887) := "00000000";
		var_ram(888) := "00000000";
		var_ram(889) := "00000000";
		var_ram(890) := "00000000";
		var_ram(891) := "00000000";
		var_ram(892) := "00000000";
		var_ram(893) := "00000000";
		var_ram(894) := "00000000";
		var_ram(895) := "00000000";
		var_ram(896) := "00000000";
		var_ram(897) := "00000000";
		var_ram(898) := "00000000";
		var_ram(899) := "00000000";
		var_ram(900) := "00000000";
		var_ram(901) := "00000000";
		var_ram(902) := "00000000";
		var_ram(903) := "00000000";
		var_ram(904) := "00000000";
		var_ram(905) := "00000000";
		var_ram(906) := "00000000";
		var_ram(907) := "00000000";
		var_ram(908) := "00000000";
		var_ram(909) := "00000000";
		var_ram(910) := "00000000";
		var_ram(911) := "00000000";
		var_ram(912) := "00000000";
		var_ram(913) := "00000000";
		var_ram(914) := "00000000";
		var_ram(915) := "00000000";
		var_ram(916) := "00000000";
		var_ram(917) := "00000000";
		var_ram(918) := "00000000";
		var_ram(919) := "00000000";
		var_ram(920) := "00000000";
		var_ram(921) := "00000000";
		var_ram(922) := "00000000";
		var_ram(923) := "00000000";
		var_ram(924) := "00000000";
		var_ram(925) := "00000000";
		var_ram(926) := "00000000";
		var_ram(927) := "00000000";
		var_ram(928) := "00000000";
		var_ram(929) := "00000000";
		var_ram(930) := "00000000";
		var_ram(931) := "00000000";
		var_ram(932) := "00000000";
		var_ram(933) := "00000000";
		var_ram(934) := "00000000";
		var_ram(935) := "00000000";
		var_ram(936) := "00000000";
		var_ram(937) := "00000000";
		var_ram(938) := "00000000";
		var_ram(939) := "00000000";
		var_ram(940) := "00000000";
		var_ram(941) := "00000000";
		var_ram(942) := "00000000";
		var_ram(943) := "00000000";
		var_ram(944) := "00000000";
		var_ram(945) := "00000000";
		var_ram(946) := "00000000";
		var_ram(947) := "00000000";
		var_ram(948) := "00000000";
		var_ram(949) := "00000000";
		var_ram(950) := "00000000";
		var_ram(951) := "00000000";
		var_ram(952) := "00000000";
		var_ram(953) := "00000000";
		var_ram(954) := "00000000";
		var_ram(955) := "00000000";
		var_ram(956) := "00000000";
		var_ram(957) := "00000000";
		var_ram(958) := "00000000";
		var_ram(959) := "00000000";
		var_ram(960) := "00000000";
		var_ram(961) := "00000000";
		var_ram(962) := "00000000";
		var_ram(963) := "00000000";
		var_ram(964) := "00000000";
		var_ram(965) := "00000000";
		var_ram(966) := "00000000";
		var_ram(967) := "00000000";
		var_ram(968) := "00000000";
		var_ram(969) := "00000000";
		var_ram(970) := "00000000";
		var_ram(971) := "00000000";
		var_ram(972) := "00000000";
		var_ram(973) := "00000000";
		var_ram(974) := "00000000";
		var_ram(975) := "00000000";
		var_ram(976) := "00000000";
		var_ram(977) := "00000000";
		var_ram(978) := "00000000";
		var_ram(979) := "00000000";
		var_ram(980) := "00000000";
		var_ram(981) := "00000000";
		var_ram(982) := "00000000";
		var_ram(983) := "00000000";
		var_ram(984) := "00000000";
		var_ram(985) := "00000000";
		var_ram(986) := "00000000";
		var_ram(987) := "00000000";
		var_ram(988) := "00000000";
		var_ram(989) := "00000000";
		var_ram(990) := "00000000";
		var_ram(991) := "00000000";
		var_ram(992) := "00000000";
		var_ram(993) := "00000000";
		var_ram(994) := "00000000";
		var_ram(995) := "00000000";
		var_ram(996) := "00000000";
		var_ram(997) := "00000000";
		var_ram(998) := "00000000";
		var_ram(999) := "00000000";
		var_ram(1000) := "00000000";
		var_ram(1001) := "00000000";
		var_ram(1002) := "00000000";
		var_ram(1003) := "00000000";
		var_ram(1004) := "00000000";
		var_ram(1005) := "00000000";
		var_ram(1006) := "00000000";
		var_ram(1007) := "00000000";
		var_ram(1008) := "00000000";
		var_ram(1009) := "00000000";
		var_ram(1010) := "00000000";
		var_ram(1011) := "00000000";
		var_ram(1012) := "00000000";
		var_ram(1013) := "00000000";
		var_ram(1014) := "00000000";
		var_ram(1015) := "00000000";
		var_ram(1016) := "00000000";
		var_ram(1017) := "00000000";
		var_ram(1018) := "00000000";
		var_ram(1019) := "00000000";
		var_ram(1020) := "00000000";
		var_ram(1021) := "00000000";
		var_ram(1022) := "00000000";
		var_ram(1023) := "00000000";
		var_ram(1024) := "00000000";
		var_ram(1025) := "00000000";
		var_ram(1026) := "00000000";
		var_ram(1027) := "00000000";
		var_ram(1028) := "00000000";
		var_ram(1029) := "00000000";
		var_ram(1030) := "00000000";
		var_ram(1031) := "00000000";
		var_ram(1032) := "00000000";
		var_ram(1033) := "00000000";
		var_ram(1034) := "00000000";
		var_ram(1035) := "00000000";
		var_ram(1036) := "00000000";
		var_ram(1037) := "00000000";
		var_ram(1038) := "00000000";
		var_ram(1039) := "00000000";
		var_ram(1040) := "00000000";
		var_ram(1041) := "00000000";
		var_ram(1042) := "00000000";
		var_ram(1043) := "00000000";
		var_ram(1044) := "00000000";
		var_ram(1045) := "00000000";
		var_ram(1046) := "00000000";
		var_ram(1047) := "00000000";
		var_ram(1048) := "00000000";
		var_ram(1049) := "00000000";
		var_ram(1050) := "00000000";
		var_ram(1051) := "00000000";
		var_ram(1052) := "00000000";
		var_ram(1053) := "00000000";
		var_ram(1054) := "00000000";
		var_ram(1055) := "00000000";
		var_ram(1056) := "00000000";
		var_ram(1057) := "00000000";
		var_ram(1058) := "00000000";
		var_ram(1059) := "00000000";
		var_ram(1060) := "00000000";
		var_ram(1061) := "00000000";
		var_ram(1062) := "00000000";
		var_ram(1063) := "00000000";
		var_ram(1064) := "00000000";
		var_ram(1065) := "00000000";
		var_ram(1066) := "00000000";
		var_ram(1067) := "00000000";
		var_ram(1068) := "00000000";
		var_ram(1069) := "00000000";
		var_ram(1070) := "00000000";
		var_ram(1071) := "00000000";
		var_ram(1072) := "00000000";
		var_ram(1073) := "00000000";
		var_ram(1074) := "00000000";
		var_ram(1075) := "00000000";
		var_ram(1076) := "00000000";
		var_ram(1077) := "00000000";
		var_ram(1078) := "00000000";
		var_ram(1079) := "00000000";
		var_ram(1080) := "00000000";
		var_ram(1081) := "00000000";
		var_ram(1082) := "00000000";
		var_ram(1083) := "00000000";
		var_ram(1084) := "00000000";
		var_ram(1085) := "00000000";
		var_ram(1086) := "00000000";
		var_ram(1087) := "00000000";
		var_ram(1088) := "00000000";
		var_ram(1089) := "00000000";
		var_ram(1090) := "00000000";
		var_ram(1091) := "00000000";
		var_ram(1092) := "00000000";
		var_ram(1093) := "00000000";
		var_ram(1094) := "00000000";
		var_ram(1095) := "00000000";
		var_ram(1096) := "00000000";
		var_ram(1097) := "00000000";
		var_ram(1098) := "00000000";
		var_ram(1099) := "00000000";
		var_ram(1100) := "00000000";
		var_ram(1101) := "00000000";
		var_ram(1102) := "00000000";
		var_ram(1103) := "00000000";
		var_ram(1104) := "00000000";
		var_ram(1105) := "00000000";
		var_ram(1106) := "00000000";
		var_ram(1107) := "00000000";
		var_ram(1108) := "00000000";
		var_ram(1109) := "00000000";
		var_ram(1110) := "00000000";
		var_ram(1111) := "00000000";
		var_ram(1112) := "00000000";
		var_ram(1113) := "00000000";
		var_ram(1114) := "00000000";
		var_ram(1115) := "00000000";
		var_ram(1116) := "00000000";
		var_ram(1117) := "00000000";
		var_ram(1118) := "00000000";
		var_ram(1119) := "00000000";
		var_ram(1120) := "00000000";
		var_ram(1121) := "00000000";
		var_ram(1122) := "00000000";
		var_ram(1123) := "00000000";
		var_ram(1124) := "00000000";
		var_ram(1125) := "00000000";
		var_ram(1126) := "00000000";
		var_ram(1127) := "00000000";
		var_ram(1128) := "00000000";
		var_ram(1129) := "00000000";
		var_ram(1130) := "00000000";
		var_ram(1131) := "00000000";
		var_ram(1132) := "00000000";
		var_ram(1133) := "00000000";
		var_ram(1134) := "00000000";
		var_ram(1135) := "00000000";
		var_ram(1136) := "00000000";
		var_ram(1137) := "00000000";
		var_ram(1138) := "00000000";
		var_ram(1139) := "00000000";
		var_ram(1140) := "00000000";
		var_ram(1141) := "00000000";
		var_ram(1142) := "00000000";
		var_ram(1143) := "00000000";
		var_ram(1144) := "00000000";
		var_ram(1145) := "00000000";
		var_ram(1146) := "00000000";
		var_ram(1147) := "00000000";
		var_ram(1148) := "00000000";
		var_ram(1149) := "00000000";
		var_ram(1150) := "00000000";
		var_ram(1151) := "00000000";
		var_ram(1152) := "00000000";
		var_ram(1153) := "00000000";
		var_ram(1154) := "00000000";
		var_ram(1155) := "00000000";
		var_ram(1156) := "00000000";
		var_ram(1157) := "00000000";
		var_ram(1158) := "00000000";
		var_ram(1159) := "00000000";
		var_ram(1160) := "00000000";
		var_ram(1161) := "00000000";
		var_ram(1162) := "00000000";
		var_ram(1163) := "00000000";
		var_ram(1164) := "00000000";
		var_ram(1165) := "00000000";
		var_ram(1166) := "00000000";
		var_ram(1167) := "00000000";
		var_ram(1168) := "00000000";
		var_ram(1169) := "00000000";
		var_ram(1170) := "00000000";
		var_ram(1171) := "00000000";
		var_ram(1172) := "00000000";
		var_ram(1173) := "00000000";
		var_ram(1174) := "00000000";
		var_ram(1175) := "00000000";
		var_ram(1176) := "00000000";
		var_ram(1177) := "00000000";
		var_ram(1178) := "00000000";
		var_ram(1179) := "00000000";
		var_ram(1180) := "00000000";
		var_ram(1181) := "00000000";
		var_ram(1182) := "00000000";
		var_ram(1183) := "00000000";
		var_ram(1184) := "00000000";
		var_ram(1185) := "00000000";
		var_ram(1186) := "00000000";
		var_ram(1187) := "00000000";
		var_ram(1188) := "00000000";
		var_ram(1189) := "00000000";
		var_ram(1190) := "00000000";
		var_ram(1191) := "00000000";
		var_ram(1192) := "00000000";
		var_ram(1193) := "00000000";
		var_ram(1194) := "00000000";
		var_ram(1195) := "00000000";
		var_ram(1196) := "00000000";
		var_ram(1197) := "00000000";
		var_ram(1198) := "00000000";
		var_ram(1199) := "00000000";
		var_ram(1200) := "00000000";
		var_ram(1201) := "00000000";
		var_ram(1202) := "00000000";
		var_ram(1203) := "00000000";
		var_ram(1204) := "00000000";
		var_ram(1205) := "00000000";
		var_ram(1206) := "00000000";
		var_ram(1207) := "00000000";
		var_ram(1208) := "00000000";
		var_ram(1209) := "00000000";
		var_ram(1210) := "00000000";
		var_ram(1211) := "00000000";
		var_ram(1212) := "00000000";
		var_ram(1213) := "00000000";
		var_ram(1214) := "00000000";
		var_ram(1215) := "00000000";
		var_ram(1216) := "00000000";
		var_ram(1217) := "00000000";
		var_ram(1218) := "00000000";
		var_ram(1219) := "00000000";
		var_ram(1220) := "00000000";
		var_ram(1221) := "00000000";
		var_ram(1222) := "00000000";
		var_ram(1223) := "00000000";
		var_ram(1224) := "00000000";
		var_ram(1225) := "00000000";
		var_ram(1226) := "00000000";
		var_ram(1227) := "00000000";
		var_ram(1228) := "00000000";
		var_ram(1229) := "00000000";
		var_ram(1230) := "00000000";
		var_ram(1231) := "00000000";
		var_ram(1232) := "00000000";
		var_ram(1233) := "00000000";
		var_ram(1234) := "00000000";
		var_ram(1235) := "00000000";
		var_ram(1236) := "00000000";
		var_ram(1237) := "00000000";
		var_ram(1238) := "00000000";
		var_ram(1239) := "00000000";
		var_ram(1240) := "00000000";
		var_ram(1241) := "00000000";
		var_ram(1242) := "00000000";
		var_ram(1243) := "00000000";
		var_ram(1244) := "00000000";
		var_ram(1245) := "00000000";
		var_ram(1246) := "00000000";
		var_ram(1247) := "00000000";
		var_ram(1248) := "00000000";
		var_ram(1249) := "00000000";
		var_ram(1250) := "00000000";
		var_ram(1251) := "00000000";
		var_ram(1252) := "00000000";
		var_ram(1253) := "00000000";
		var_ram(1254) := "00000000";
		var_ram(1255) := "00000000";
		var_ram(1256) := "00000000";
		var_ram(1257) := "00000000";
		var_ram(1258) := "00000000";
		var_ram(1259) := "00000000";
		var_ram(1260) := "00000000";
		var_ram(1261) := "00000000";
		var_ram(1262) := "00000000";
		var_ram(1263) := "00000000";
		var_ram(1264) := "00000000";
		var_ram(1265) := "00000000";
		var_ram(1266) := "00000000";
		var_ram(1267) := "00000000";
		var_ram(1268) := "00000000";
		var_ram(1269) := "00000000";
		var_ram(1270) := "00000000";
		var_ram(1271) := "00000000";
		var_ram(1272) := "00000000";
		var_ram(1273) := "00000000";
		var_ram(1274) := "00000000";
		var_ram(1275) := "00000000";
		var_ram(1276) := "00000000";
		var_ram(1277) := "00000000";
		var_ram(1278) := "00000000";
		var_ram(1279) := "00000000";
		var_ram(1280) := "00000000";
		var_ram(1281) := "00000000";
		var_ram(1282) := "00000000";
		var_ram(1283) := "00000000";
		var_ram(1284) := "00000000";
		var_ram(1285) := "00000000";
		var_ram(1286) := "00000000";
		var_ram(1287) := "00000000";
		var_ram(1288) := "00000000";
		var_ram(1289) := "00000000";
		var_ram(1290) := "00000000";
		var_ram(1291) := "00000000";
		var_ram(1292) := "00000000";
		var_ram(1293) := "00000000";
		var_ram(1294) := "00000000";
		var_ram(1295) := "00000000";
		var_ram(1296) := "00000000";
		var_ram(1297) := "00000000";
		var_ram(1298) := "00000000";
		var_ram(1299) := "00000000";
		var_ram(1300) := "00000000";
		var_ram(1301) := "00000000";
		var_ram(1302) := "00000000";
		var_ram(1303) := "00000000";
		var_ram(1304) := "00000000";
		var_ram(1305) := "00000000";
		var_ram(1306) := "00000000";
		var_ram(1307) := "00000000";
		var_ram(1308) := "00000000";
		var_ram(1309) := "00000000";
		var_ram(1310) := "00000000";
		var_ram(1311) := "00000000";
		var_ram(1312) := "00000000";
		var_ram(1313) := "00000000";
		var_ram(1314) := "00000000";
		var_ram(1315) := "00000000";
		var_ram(1316) := "00000000";
		var_ram(1317) := "00000000";
		var_ram(1318) := "00000000";
		var_ram(1319) := "00000000";
		var_ram(1320) := "00000000";
		var_ram(1321) := "00000000";
		var_ram(1322) := "00000000";
		var_ram(1323) := "00000000";
		var_ram(1324) := "00000000";
		var_ram(1325) := "00000000";
		var_ram(1326) := "00000000";
		var_ram(1327) := "00000000";
		var_ram(1328) := "00000000";
		var_ram(1329) := "00000000";
		var_ram(1330) := "00000000";
		var_ram(1331) := "00000000";
		var_ram(1332) := "00000000";
		var_ram(1333) := "00000000";
		var_ram(1334) := "00000000";
		var_ram(1335) := "00000000";
		var_ram(1336) := "00000000";
		var_ram(1337) := "00000000";
		var_ram(1338) := "00000000";
		var_ram(1339) := "00000000";
		var_ram(1340) := "00000000";
		var_ram(1341) := "00000000";
		var_ram(1342) := "00000000";
		var_ram(1343) := "00000000";
		var_ram(1344) := "00000000";
		var_ram(1345) := "00000000";
		var_ram(1346) := "00000000";
		var_ram(1347) := "00000000";
		var_ram(1348) := "00000000";
		var_ram(1349) := "00000000";
		var_ram(1350) := "00000000";
		var_ram(1351) := "00000000";
		var_ram(1352) := "00000000";
		var_ram(1353) := "00000000";
		var_ram(1354) := "00000000";
		var_ram(1355) := "00000000";
		var_ram(1356) := "00000000";
		var_ram(1357) := "00000000";
		var_ram(1358) := "00000000";
		var_ram(1359) := "00000000";
		var_ram(1360) := "00000000";
		var_ram(1361) := "00000000";
		var_ram(1362) := "00000000";
		var_ram(1363) := "00000000";
		var_ram(1364) := "00000000";
		var_ram(1365) := "00000000";
		var_ram(1366) := "00000000";
		var_ram(1367) := "00000000";
		var_ram(1368) := "00000000";
		var_ram(1369) := "00000000";
		var_ram(1370) := "00000000";
		var_ram(1371) := "00000000";
		var_ram(1372) := "00000000";
		var_ram(1373) := "00000000";
		var_ram(1374) := "00000000";
		var_ram(1375) := "00000000";
		var_ram(1376) := "00000000";
		var_ram(1377) := "00000000";
		var_ram(1378) := "00000000";
		var_ram(1379) := "00000000";
		var_ram(1380) := "00000000";
		var_ram(1381) := "00000000";
		var_ram(1382) := "00000000";
		var_ram(1383) := "00000000";
		var_ram(1384) := "00000000";
		var_ram(1385) := "00000000";
		var_ram(1386) := "00000000";
		var_ram(1387) := "00000000";
		var_ram(1388) := "00000000";
		var_ram(1389) := "00000000";
		var_ram(1390) := "00000000";
		var_ram(1391) := "00000000";
		var_ram(1392) := "00000000";
		var_ram(1393) := "00000000";
		var_ram(1394) := "00000000";
		var_ram(1395) := "00000000";
		var_ram(1396) := "00000000";
		var_ram(1397) := "00000000";
		var_ram(1398) := "00000000";
		var_ram(1399) := "00000000";
		var_ram(1400) := "00000000";
		var_ram(1401) := "00000000";
		var_ram(1402) := "00000000";
		var_ram(1403) := "00000000";
		var_ram(1404) := "00000000";
		var_ram(1405) := "00000000";
		var_ram(1406) := "00000000";
		var_ram(1407) := "00000000";
		var_ram(1408) := "00000000";
		var_ram(1409) := "00000000";
		var_ram(1410) := "00000000";
		var_ram(1411) := "00000000";
		var_ram(1412) := "00000000";
		var_ram(1413) := "00000000";
		var_ram(1414) := "00000000";
		var_ram(1415) := "00000000";
		var_ram(1416) := "00000000";
		var_ram(1417) := "00000000";
		var_ram(1418) := "00000000";
		var_ram(1419) := "00000000";
		var_ram(1420) := "00000000";
		var_ram(1421) := "00000000";
		var_ram(1422) := "00000000";
		var_ram(1423) := "00000000";
		var_ram(1424) := "00000000";
		var_ram(1425) := "00000000";
		var_ram(1426) := "00000000";
		var_ram(1427) := "00000000";
		var_ram(1428) := "00000000";
		var_ram(1429) := "00000000";
		var_ram(1430) := "00000000";
		var_ram(1431) := "00000000";
		var_ram(1432) := "00000000";
		var_ram(1433) := "00000000";
		var_ram(1434) := "00000000";
		var_ram(1435) := "00000000";
		var_ram(1436) := "00000000";
		var_ram(1437) := "00000000";
		var_ram(1438) := "00000000";
		var_ram(1439) := "00000000";
		var_ram(1440) := "00000000";
		var_ram(1441) := "00000000";
		var_ram(1442) := "00000000";
		var_ram(1443) := "00000000";
		var_ram(1444) := "00000000";
		var_ram(1445) := "00000000";
		var_ram(1446) := "00000000";
		var_ram(1447) := "00000000";
		var_ram(1448) := "00000000";
		var_ram(1449) := "00000000";
		var_ram(1450) := "00000000";
		var_ram(1451) := "00000000";
		var_ram(1452) := "00000000";
		var_ram(1453) := "00000000";
		var_ram(1454) := "00000000";
		var_ram(1455) := "00000000";
		var_ram(1456) := "00000000";
		var_ram(1457) := "00000000";
		var_ram(1458) := "00000000";
		var_ram(1459) := "00000000";
		var_ram(1460) := "00000000";
		var_ram(1461) := "00000000";
		var_ram(1462) := "00000000";
		var_ram(1463) := "00000000";
		var_ram(1464) := "00000000";
		var_ram(1465) := "00000000";
		var_ram(1466) := "00000000";
		var_ram(1467) := "00000000";
		var_ram(1468) := "00000000";
		var_ram(1469) := "00000000";
		var_ram(1470) := "00000000";
		var_ram(1471) := "00000000";
		var_ram(1472) := "00000000";
		var_ram(1473) := "00000000";
		var_ram(1474) := "00000000";
		var_ram(1475) := "00000000";
		var_ram(1476) := "00000000";
		var_ram(1477) := "00000000";
		var_ram(1478) := "00000000";
		var_ram(1479) := "00000000";
		var_ram(1480) := "00000000";
		var_ram(1481) := "00000000";
		var_ram(1482) := "00000000";
		var_ram(1483) := "00000000";
		var_ram(1484) := "00000000";
		var_ram(1485) := "00000000";
		var_ram(1486) := "00000000";
		var_ram(1487) := "00000000";
		var_ram(1488) := "00000000";
		var_ram(1489) := "00000000";
		var_ram(1490) := "00000000";
		var_ram(1491) := "00000000";
		var_ram(1492) := "00000000";
		var_ram(1493) := "00000000";
		var_ram(1494) := "00000000";
		var_ram(1495) := "00000000";
		var_ram(1496) := "00000000";
		var_ram(1497) := "00000000";
		var_ram(1498) := "00000000";
		var_ram(1499) := "00000000";
		var_ram(1500) := "00000000";
		var_ram(1501) := "00000000";
		var_ram(1502) := "00000000";
		var_ram(1503) := "00000000";
		var_ram(1504) := "00000000";
		var_ram(1505) := "00000000";
		var_ram(1506) := "00000000";
		var_ram(1507) := "00000000";
		var_ram(1508) := "00000000";
		var_ram(1509) := "00000000";
		var_ram(1510) := "00000000";
		var_ram(1511) := "00000000";
		var_ram(1512) := "00000000";
		var_ram(1513) := "00000000";
		var_ram(1514) := "00000000";
		var_ram(1515) := "00000000";
		var_ram(1516) := "00000000";
		var_ram(1517) := "00000000";
		var_ram(1518) := "00000000";
		var_ram(1519) := "00000000";
		var_ram(1520) := "00000000";
		var_ram(1521) := "00000000";
		var_ram(1522) := "00000000";
		var_ram(1523) := "00000000";
		var_ram(1524) := "00000000";
		var_ram(1525) := "00000000";
		var_ram(1526) := "00000000";
		var_ram(1527) := "00000000";
		var_ram(1528) := "00000000";
		var_ram(1529) := "00000000";
		var_ram(1530) := "00000000";
		var_ram(1531) := "00000000";
		var_ram(1532) := "00000000";
		var_ram(1533) := "00000000";
		var_ram(1534) := "00000000";
		var_ram(1535) := "00000000";
		var_ram(1536) := "00000000";
		var_ram(1537) := "00000000";
		var_ram(1538) := "00000000";
		var_ram(1539) := "00000000";
		var_ram(1540) := "00000000";
		var_ram(1541) := "00000000";
		var_ram(1542) := "00000000";
		var_ram(1543) := "00000000";
		var_ram(1544) := "00000000";
		var_ram(1545) := "00000000";
		var_ram(1546) := "00000000";
		var_ram(1547) := "00000000";
		var_ram(1548) := "00000000";
		var_ram(1549) := "00000000";
		var_ram(1550) := "00000000";
		var_ram(1551) := "00000000";
		var_ram(1552) := "00000000";
		var_ram(1553) := "00000000";
		var_ram(1554) := "00000000";
		var_ram(1555) := "00000000";
		var_ram(1556) := "00000000";
		var_ram(1557) := "00000000";
		var_ram(1558) := "00000000";
		var_ram(1559) := "00000000";
		var_ram(1560) := "00000000";
		var_ram(1561) := "00000000";
		var_ram(1562) := "00000000";
		var_ram(1563) := "00000000";
		var_ram(1564) := "00000000";
		var_ram(1565) := "00000000";
		var_ram(1566) := "00000000";
		var_ram(1567) := "00000000";
		var_ram(1568) := "00000000";
		var_ram(1569) := "00000000";
		var_ram(1570) := "00000000";
		var_ram(1571) := "00000000";
		var_ram(1572) := "00000000";
		var_ram(1573) := "00000000";
		var_ram(1574) := "00000000";
		var_ram(1575) := "00000000";
		var_ram(1576) := "00000000";
		var_ram(1577) := "00000000";
		var_ram(1578) := "00000000";
		var_ram(1579) := "00000000";
		var_ram(1580) := "00000000";
		var_ram(1581) := "00000000";
		var_ram(1582) := "00000000";
		var_ram(1583) := "00000000";
		var_ram(1584) := "00000000";
		var_ram(1585) := "00000000";
		var_ram(1586) := "00000000";
		var_ram(1587) := "00000000";
		var_ram(1588) := "00000000";
		var_ram(1589) := "00000000";
		var_ram(1590) := "00000000";
		var_ram(1591) := "00000000";
		var_ram(1592) := "00000000";
		var_ram(1593) := "00000000";
		var_ram(1594) := "00000000";
		var_ram(1595) := "00000000";
		var_ram(1596) := "00000000";
		var_ram(1597) := "00000000";
		var_ram(1598) := "00000000";
		var_ram(1599) := "00000000";
		var_ram(1600) := "00000000";
		var_ram(1601) := "00000000";
		var_ram(1602) := "00000000";
		var_ram(1603) := "00000000";
		var_ram(1604) := "00000000";
		var_ram(1605) := "00000000";
		var_ram(1606) := "00000000";
		var_ram(1607) := "00000000";
		var_ram(1608) := "00000000";
		var_ram(1609) := "00000000";
		var_ram(1610) := "00000000";
		var_ram(1611) := "00000000";
		var_ram(1612) := "00000000";
		var_ram(1613) := "00000000";
		var_ram(1614) := "00000000";
		var_ram(1615) := "00000000";
		var_ram(1616) := "00000000";
		var_ram(1617) := "00000000";
		var_ram(1618) := "00000000";
		var_ram(1619) := "00000000";
		var_ram(1620) := "00000000";
		var_ram(1621) := "00000000";
		var_ram(1622) := "00000000";
		var_ram(1623) := "00000000";
		var_ram(1624) := "00000000";
		var_ram(1625) := "00000000";
		var_ram(1626) := "00000000";
		var_ram(1627) := "00000000";
		var_ram(1628) := "00000000";
		var_ram(1629) := "00000000";
		var_ram(1630) := "00000000";
		var_ram(1631) := "00000000";
		var_ram(1632) := "00000000";
		var_ram(1633) := "00000000";
		var_ram(1634) := "00000000";
		var_ram(1635) := "00000000";
		var_ram(1636) := "00000000";
		var_ram(1637) := "00000000";
		var_ram(1638) := "00000000";
		var_ram(1639) := "00000000";
		var_ram(1640) := "00000000";
		var_ram(1641) := "00000000";
		var_ram(1642) := "00000000";
		var_ram(1643) := "00000000";
		var_ram(1644) := "00000000";
		var_ram(1645) := "00000000";
		var_ram(1646) := "00000000";
		var_ram(1647) := "00000000";
		var_ram(1648) := "00000000";
		var_ram(1649) := "00000000";
		var_ram(1650) := "00000000";
		var_ram(1651) := "00000000";
		var_ram(1652) := "00000000";
		var_ram(1653) := "00000000";
		var_ram(1654) := "00000000";
		var_ram(1655) := "00000000";
		var_ram(1656) := "00000000";
		var_ram(1657) := "00000000";
		var_ram(1658) := "00000000";
		var_ram(1659) := "00000000";
		var_ram(1660) := "00000000";
		var_ram(1661) := "00000000";
		var_ram(1662) := "00000000";
		var_ram(1663) := "00000000";
		var_ram(1664) := "00000000";
		var_ram(1665) := "00000000";
		var_ram(1666) := "00000000";
		var_ram(1667) := "00000000";
		var_ram(1668) := "00000000";
		var_ram(1669) := "00000000";
		var_ram(1670) := "00000000";
		var_ram(1671) := "00000000";
		var_ram(1672) := "00000000";
		var_ram(1673) := "00000000";
		var_ram(1674) := "00000000";
		var_ram(1675) := "00000000";
		var_ram(1676) := "00000000";
		var_ram(1677) := "00000000";
		var_ram(1678) := "00000000";
		var_ram(1679) := "00000000";
		var_ram(1680) := "00000000";
		var_ram(1681) := "00000000";
		var_ram(1682) := "00000000";
		var_ram(1683) := "00000000";
		var_ram(1684) := "00000000";
		var_ram(1685) := "00000000";
		var_ram(1686) := "00000000";
		var_ram(1687) := "00000000";
		var_ram(1688) := "00000000";
		var_ram(1689) := "00000000";
		var_ram(1690) := "00000000";
		var_ram(1691) := "00000000";
		var_ram(1692) := "00000000";
		var_ram(1693) := "00000000";
		var_ram(1694) := "00000000";
		var_ram(1695) := "00000000";
		var_ram(1696) := "00000000";
		var_ram(1697) := "00000000";
		var_ram(1698) := "00000000";
		var_ram(1699) := "00000000";
		var_ram(1700) := "00000000";
		var_ram(1701) := "00000000";
		var_ram(1702) := "00000000";
		var_ram(1703) := "00000000";
		var_ram(1704) := "00000000";
		var_ram(1705) := "00000000";
		var_ram(1706) := "00000000";
		var_ram(1707) := "00000000";
		var_ram(1708) := "00000000";
		var_ram(1709) := "00000000";
		var_ram(1710) := "00000000";
		var_ram(1711) := "00000000";
		var_ram(1712) := "00000000";
		var_ram(1713) := "00000000";
		var_ram(1714) := "00000000";
		var_ram(1715) := "00000000";
		var_ram(1716) := "00000000";
		var_ram(1717) := "00000000";
		var_ram(1718) := "00000000";
		var_ram(1719) := "00000000";
		var_ram(1720) := "00000000";
		var_ram(1721) := "00000000";
		var_ram(1722) := "00000000";
		var_ram(1723) := "00000000";
		var_ram(1724) := "00000000";
		var_ram(1725) := "00000000";
		var_ram(1726) := "00000000";
		var_ram(1727) := "00000000";
		var_ram(1728) := "00000000";
		var_ram(1729) := "00000000";
		var_ram(1730) := "00000000";
		var_ram(1731) := "00000000";
		var_ram(1732) := "00000000";
		var_ram(1733) := "00000000";
		var_ram(1734) := "00000000";
		var_ram(1735) := "00000000";
		var_ram(1736) := "00000000";
		var_ram(1737) := "00000000";
		var_ram(1738) := "00000000";
		var_ram(1739) := "00000000";
		var_ram(1740) := "00000000";
		var_ram(1741) := "00000000";
		var_ram(1742) := "00000000";
		var_ram(1743) := "00000000";
		var_ram(1744) := "00000000";
		var_ram(1745) := "00000000";
		var_ram(1746) := "00000000";
		var_ram(1747) := "00000000";
		var_ram(1748) := "00000000";
		var_ram(1749) := "00000000";
		var_ram(1750) := "00000000";
		var_ram(1751) := "00000000";
		var_ram(1752) := "00000000";
		var_ram(1753) := "00000000";
		var_ram(1754) := "00000000";
		var_ram(1755) := "00000000";
		var_ram(1756) := "00000000";
		var_ram(1757) := "00000000";
		var_ram(1758) := "00000000";
		var_ram(1759) := "00000000";
		var_ram(1760) := "00000000";
		var_ram(1761) := "00000000";
		var_ram(1762) := "00000000";
		var_ram(1763) := "00000000";
		var_ram(1764) := "00000000";
		var_ram(1765) := "00000000";
		var_ram(1766) := "00000000";
		var_ram(1767) := "00000000";
		var_ram(1768) := "00000000";
		var_ram(1769) := "00000000";
		var_ram(1770) := "00000000";
		var_ram(1771) := "00000000";
		var_ram(1772) := "00000000";
		var_ram(1773) := "00000000";
		var_ram(1774) := "00000000";
		var_ram(1775) := "00000000";
		var_ram(1776) := "00000000";
		var_ram(1777) := "00000000";
		var_ram(1778) := "00000000";
		var_ram(1779) := "00000000";
		var_ram(1780) := "00000000";
		var_ram(1781) := "00000000";
		var_ram(1782) := "00000000";
		var_ram(1783) := "00000000";
		var_ram(1784) := "00000000";
		var_ram(1785) := "00000000";
		var_ram(1786) := "00000000";
		var_ram(1787) := "00000000";
		var_ram(1788) := "00000000";
		var_ram(1789) := "00000000";
		var_ram(1790) := "00000000";
		var_ram(1791) := "00000000";
		var_ram(1792) := "00000000";
		var_ram(1793) := "00000000";
		var_ram(1794) := "00000000";
		var_ram(1795) := "00000000";
		var_ram(1796) := "00000000";
		var_ram(1797) := "00000000";
		var_ram(1798) := "00000000";
		var_ram(1799) := "00000000";
		var_ram(1800) := "00000000";
		var_ram(1801) := "00000000";
		var_ram(1802) := "00000000";
		var_ram(1803) := "00000000";
		var_ram(1804) := "00000000";
		var_ram(1805) := "00000000";
		var_ram(1806) := "00000000";
		var_ram(1807) := "00000000";
		var_ram(1808) := "00000000";
		var_ram(1809) := "00000000";
		var_ram(1810) := "00000000";
		var_ram(1811) := "00000000";
		var_ram(1812) := "00000000";
		var_ram(1813) := "00000000";
		var_ram(1814) := "00000000";
		var_ram(1815) := "00000000";
		var_ram(1816) := "00000000";
		var_ram(1817) := "00000000";
		var_ram(1818) := "00000000";
		var_ram(1819) := "00000000";
		var_ram(1820) := "00000000";
		var_ram(1821) := "00000000";
		var_ram(1822) := "00000000";
		var_ram(1823) := "00000000";
		var_ram(1824) := "00000000";
		var_ram(1825) := "00000000";
		var_ram(1826) := "00000000";
		var_ram(1827) := "00000000";
		var_ram(1828) := "00000000";
		var_ram(1829) := "00000000";
		var_ram(1830) := "00000000";
		var_ram(1831) := "00000000";
		var_ram(1832) := "00000000";
		var_ram(1833) := "00000000";
		var_ram(1834) := "00000000";
		var_ram(1835) := "00000000";
		var_ram(1836) := "00000000";
		var_ram(1837) := "00000000";
		var_ram(1838) := "00000000";
		var_ram(1839) := "00000000";
		var_ram(1840) := "00000000";
		var_ram(1841) := "00000000";
		var_ram(1842) := "00000000";
		var_ram(1843) := "00000000";
		var_ram(1844) := "00000000";
		var_ram(1845) := "00000000";
		var_ram(1846) := "00000000";
		var_ram(1847) := "00000000";
		var_ram(1848) := "00000000";
		var_ram(1849) := "00000000";
		var_ram(1850) := "00000000";
		var_ram(1851) := "00000000";
		var_ram(1852) := "00000000";
		var_ram(1853) := "00000000";
		var_ram(1854) := "00000000";
		var_ram(1855) := "00000000";
		var_ram(1856) := "00000000";
		var_ram(1857) := "00000000";
		var_ram(1858) := "00000000";
		var_ram(1859) := "00000000";
		var_ram(1860) := "00000000";
		var_ram(1861) := "00000000";
		var_ram(1862) := "00000000";
		var_ram(1863) := "00000000";
		var_ram(1864) := "00000000";
		var_ram(1865) := "00000000";
		var_ram(1866) := "00000000";
		var_ram(1867) := "00000000";
		var_ram(1868) := "00000000";
		var_ram(1869) := "00000000";
		var_ram(1870) := "00000000";
		var_ram(1871) := "00000000";
		var_ram(1872) := "00000000";
		var_ram(1873) := "00000000";
		var_ram(1874) := "00000000";
		var_ram(1875) := "00000000";
		var_ram(1876) := "00000000";
		var_ram(1877) := "00000000";
		var_ram(1878) := "00000000";
		var_ram(1879) := "00000000";
		var_ram(1880) := "00000000";
		var_ram(1881) := "00000000";
		var_ram(1882) := "00000000";
		var_ram(1883) := "00000000";
		var_ram(1884) := "00000000";
		var_ram(1885) := "00000000";
		var_ram(1886) := "00000000";
		var_ram(1887) := "00000000";
		var_ram(1888) := "00000000";
		var_ram(1889) := "00000000";
		var_ram(1890) := "00000000";
		var_ram(1891) := "00000000";
		var_ram(1892) := "00000000";
		var_ram(1893) := "00000000";
		var_ram(1894) := "00000000";
		var_ram(1895) := "00000000";
		var_ram(1896) := "00000000";
		var_ram(1897) := "00000000";
		var_ram(1898) := "00000000";
		var_ram(1899) := "00000000";
		var_ram(1900) := "00000000";
		var_ram(1901) := "00000000";
		var_ram(1902) := "00000000";
		var_ram(1903) := "00000000";
		var_ram(1904) := "00000000";
		var_ram(1905) := "00000000";
		var_ram(1906) := "00000000";
		var_ram(1907) := "00000000";
		var_ram(1908) := "00000000";
		var_ram(1909) := "00000000";
		var_ram(1910) := "00000000";
		var_ram(1911) := "00000000";
		var_ram(1912) := "00000000";
		var_ram(1913) := "00000000";
		var_ram(1914) := "00000000";
		var_ram(1915) := "00000000";
		var_ram(1916) := "00000000";
		var_ram(1917) := "00000000";
		var_ram(1918) := "00000000";
		var_ram(1919) := "00000000";
		var_ram(1920) := "00000000";
		var_ram(1921) := "00000000";
		var_ram(1922) := "00000000";
		var_ram(1923) := "00000000";
		var_ram(1924) := "00000000";
		var_ram(1925) := "00000000";
		var_ram(1926) := "00000000";
		var_ram(1927) := "00000000";
		var_ram(1928) := "00000000";
		var_ram(1929) := "00000000";
		var_ram(1930) := "00000000";
		var_ram(1931) := "00000000";
		var_ram(1932) := "00000000";
		var_ram(1933) := "00000000";
		var_ram(1934) := "00000000";
		var_ram(1935) := "00000000";
		var_ram(1936) := "00000000";
		var_ram(1937) := "00000000";
		var_ram(1938) := "00000000";
		var_ram(1939) := "00000000";
		var_ram(1940) := "00000000";
		var_ram(1941) := "00000000";
		var_ram(1942) := "00000000";
		var_ram(1943) := "00000000";
		var_ram(1944) := "00000000";
		var_ram(1945) := "00000000";
		var_ram(1946) := "00000000";
		var_ram(1947) := "00000000";
		var_ram(1948) := "00000000";
		var_ram(1949) := "00000000";
		var_ram(1950) := "00000000";
		var_ram(1951) := "00000000";
		var_ram(1952) := "00000000";
		var_ram(1953) := "00000000";
		var_ram(1954) := "00000000";
		var_ram(1955) := "00000000";
		var_ram(1956) := "00000000";
		var_ram(1957) := "00000000";
		var_ram(1958) := "00000000";
		var_ram(1959) := "00000000";
		var_ram(1960) := "00000000";
		var_ram(1961) := "00000000";
		var_ram(1962) := "00000000";
		var_ram(1963) := "00000000";
		var_ram(1964) := "00000000";
		var_ram(1965) := "00000000";
		var_ram(1966) := "00000000";
		var_ram(1967) := "00000000";
		var_ram(1968) := "00000000";
		var_ram(1969) := "00000000";
		var_ram(1970) := "00000000";
		var_ram(1971) := "00000000";
		var_ram(1972) := "00000000";
		var_ram(1973) := "00000000";
		var_ram(1974) := "00000000";
		var_ram(1975) := "00000000";
		var_ram(1976) := "00000000";
		var_ram(1977) := "00000000";
		var_ram(1978) := "00000000";
		var_ram(1979) := "00000000";
		var_ram(1980) := "00000000";
		var_ram(1981) := "00000000";
		var_ram(1982) := "00000000";
		var_ram(1983) := "00000000";
		var_ram(1984) := "00000000";
		var_ram(1985) := "00000000";
		var_ram(1986) := "00000000";
		var_ram(1987) := "00000000";
		var_ram(1988) := "00000000";
		var_ram(1989) := "00000000";
		var_ram(1990) := "00000000";
		var_ram(1991) := "00000000";
		var_ram(1992) := "00000000";
		var_ram(1993) := "00000000";
		var_ram(1994) := "00000000";
		var_ram(1995) := "00000000";
		var_ram(1996) := "00000000";
		var_ram(1997) := "00000000";
		var_ram(1998) := "00000000";
		var_ram(1999) := "00000000";
		var_ram(2000) := "00000000";
		var_ram(2001) := "00000000";
		var_ram(2002) := "00000000";
		var_ram(2003) := "00000000";
		var_ram(2004) := "00000000";
		var_ram(2005) := "00000000";
		var_ram(2006) := "00000000";
		var_ram(2007) := "00000000";
		var_ram(2008) := "00000000";
		var_ram(2009) := "00000000";
		var_ram(2010) := "00000000";
		var_ram(2011) := "00000000";
		var_ram(2012) := "00000000";
		var_ram(2013) := "00000000";
		var_ram(2014) := "00000000";
		var_ram(2015) := "00000000";
		var_ram(2016) := "00000000";
		var_ram(2017) := "00000000";
		var_ram(2018) := "00000000";
		var_ram(2019) := "00000000";
		var_ram(2020) := "00000000";
		var_ram(2021) := "00000000";
		var_ram(2022) := "00000000";
		var_ram(2023) := "00000000";
		var_ram(2024) := "00000000";
		var_ram(2025) := "00000000";
		var_ram(2026) := "00000000";
		var_ram(2027) := "00000000";
		var_ram(2028) := "00000000";
		var_ram(2029) := "00000000";
		var_ram(2030) := "00000000";
		var_ram(2031) := "00000000";
		var_ram(2032) := "00000000";
		var_ram(2033) := "00000000";
		var_ram(2034) := "00000000";
		var_ram(2035) := "00000000";
		var_ram(2036) := "00000000";
		var_ram(2037) := "00000000";
		var_ram(2038) := "00000000";
		var_ram(2039) := "00000000";
		var_ram(2040) := "00000000";
		var_ram(2041) := "00000000";
		var_ram(2042) := "00000000";
		var_ram(2043) := "00000000";
		var_ram(2044) := "00000000";
		var_ram(2045) := "00000000";
		var_ram(2046) := "00000000";
		var_ram(2047) := "00000000";

		
		elsif (falling_edge(clk)) then
			var_addr := conv_integer(addr);
			if wr_en = '1' then
				var_ram(var_addr) := data_in;
			end if;
				data_out <= var_ram(var_addr);
		end if;	
		
	
	end process;
end Behavioral;

