----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date:    14:24:35 10/08/2019 
-- Design Name: 
-- Module Name:    rom - Behavioral 
-- Project Name: 
-- Target Devices: 
-- Tool versions: 
-- Description: 
--
-- Dependencies: 
--
-- Revision: 
-- Revision 0.01 - File Created
-- Additional Comments: 
--
----------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--use IEEE.NUMERIC_STD.ALL;

-- Uncomment the following library declaration if instantiating
-- any Xilinx primitives in this code.
--library UNISIM;
--use UNISIM.VComponents.all;

--named rom but is actually ram
entity ram is
    Port ( clk : in  STD_LOGIC;
           --rst : in  STD_LOGIC;
			  wr_en : in STD_LOGIC;
           addr : in  STD_LOGIC_VECTOR (9 downto 0);
			  data_in : in STD_LOGIC_VECTOR(7 downto 0);
           data_out : out  STD_LOGIC_VECTOR (7 downto 0));
end ram;

architecture Behavioral of ram is

type ram_type is array (0 to 1023) of std_logic_vector(7 downto 0);
signal ram : ram_type := (others => (others => '0'));

begin

	ram_process: process(clk, addr) is
	--variable var_ram : ram_type;
	variable var_addr : integer;
	
	begin
--		if (rst = '1') then
--		
--			ram(0) <= "00000000";
--			ram(1) <= "00000000";
--			ram(2) <= "00000000";
--			ram(3) <= "00000000";
--			ram(4) <= "00000000";
--			ram(5) <= "00000000";
--			ram(6) <= "00000000";
--			ram(7) <= "00000000";
--			ram(8) <= "00000000";
--			ram(9) <= "00000000";
--			ram(10) <= "00000000";
--			ram(11) <= "00000000";
--			ram(12) <= "00000000";
--			ram(13) <= "00000000";
--			ram(14) <= "00000000";
--			ram(15) <= "00000000";
--			ram(16) <= "00000000";
--			ram(17) <= "00000000";
--			ram(18) <= "00000000";
--			ram(19) <= "00000000";
--			ram(20) <= "00000000";
--			ram(21) <= "00000000";
--			ram(22) <= "00000000";
--			ram(23) <= "00000000";
--			ram(24) <= "00000000";
--			ram(25) <= "00000000";
--			ram(26) <= "00000000";
--			ram(27) <= "00000000";
--			ram(28) <= "00000000";
--			ram(29) <= "00000000";
--			ram(30) <= "00000000";
--			ram(31) <= "00000000";
--			ram(32) <= "00000000";
--			ram(33) <= "00000000";
--			ram(34) <= "00000000";
--			ram(35) <= "00000000";
--			ram(36) <= "00000000";
--			ram(37) <= "00000000";
--			ram(38) <= "00000000";
--			ram(39) <= "00000000";
--			ram(40) <= "00000000";
--			ram(41) <= "00000000";
--			ram(42) <= "00000000";
--			ram(43) <= "00000000";
--			ram(44) <= "00000000";
--			ram(45) <= "00000000";
--			ram(46) <= "00000000";
--			ram(47) <= "00000000";
--			ram(48) <= "00000000";
--			ram(49) <= "00000000";
--			ram(50) <= "00000000";
--			ram(51) <= "00000000";
--			ram(52) <= "00000000";
--			ram(53) <= "00000000";
--			ram(54) <= "00000000";
--			ram(55) <= "00000000";
--			ram(56) <= "00000000";
--			ram(57) <= "00000000";
--			ram(58) <= "00000000";
--			ram(59) <= "00000000";
--			ram(60) <= "00000000";
--			ram(61) <= "00000000";
--			ram(62) <= "00000000";
--			ram(63) <= "00000000";
--			ram(64) <= "00000000";
--			ram(65) <= "00000000";
--			ram(66) <= "00000000";
--			ram(67) <= "00000000";
--			ram(68) <= "00000000";
--			ram(69) <= "00000000";
--			ram(70) <= "00000000";
--			ram(71) <= "00000000";
--			ram(72) <= "00000000";
--			ram(73) <= "00000000";
--			ram(74) <= "00000000";
--			ram(75) <= "00000000";
--			ram(76) <= "00000000";
--			ram(77) <= "00000000";
--			ram(78) <= "00000000";
--			ram(79) <= "00000000";
--			ram(80) <= "00000000";
--			ram(81) <= "00000000";
--			ram(82) <= "00000000";
--			ram(83) <= "00000000";
--			ram(84) <= "00000000";
--			ram(85) <= "00000000";
--			ram(86) <= "00000000";
--			ram(87) <= "00000000";
--			ram(88) <= "00000000";
--			ram(89) <= "00000000";
--			ram(90) <= "00000000";
--			ram(91) <= "00000000";
--			ram(92) <= "00000000";
--			ram(93) <= "00000000";
--			ram(94) <= "00000000";
--			ram(95) <= "00000000";
--			ram(96) <= "00000000";
--			ram(97) <= "00000000";
--			ram(98) <= "00000000";
--			ram(99) <= "00000000";
--			ram(100) <= "00000000";
--			ram(101) <= "00000000";
--			ram(102) <= "00000000";
--			ram(103) <= "00000000";
--			ram(104) <= "00000000";
--			ram(105) <= "00000000";
--			ram(106) <= "00000000";
--			ram(107) <= "00000000";
--			ram(108) <= "00000000";
--			ram(109) <= "00000000";
--			ram(110) <= "00000000";
--			ram(111) <= "00000000";
--			ram(112) <= "00000000";
--			ram(113) <= "00000000";
--			ram(114) <= "00000000";
--			ram(115) <= "00000000";
--			ram(116) <= "00000000";
--			ram(117) <= "00000000";
--			ram(118) <= "00000000";
--			ram(119) <= "00000000";
--			ram(120) <= "00000000";
--			ram(121) <= "00000000";
--			ram(122) <= "00000000";
--			ram(123) <= "00000000";
--			ram(124) <= "00000000";
--			ram(125) <= "00000000";
--			ram(126) <= "00000000";
--			ram(127) <= "00000000";
--			ram(128) <= "00000000";
--			ram(129) <= "00000000";
--			ram(130) <= "00000000";
--			ram(131) <= "00000000";
--			ram(132) <= "00000000";
--			ram(133) <= "00000000";
--			ram(134) <= "00000000";
--			ram(135) <= "00000000";
--			ram(136) <= "00000000";
--			ram(137) <= "00000000";
--			ram(138) <= "00000000";
--			ram(139) <= "00000000";
--			ram(140) <= "00000000";
--			ram(141) <= "00000000";
--			ram(142) <= "00000000";
--			ram(143) <= "00000000";
--			ram(144) <= "00000000";
--			ram(145) <= "00000000";
--			ram(146) <= "00000000";
--			ram(147) <= "00000000";
--			ram(148) <= "00000000";
--			ram(149) <= "00000000";
--			ram(150) <= "00000000";
--			ram(151) <= "00000000";
--			ram(152) <= "00000000";
--			ram(153) <= "00000000";
--			ram(154) <= "00000000";
--			ram(155) <= "00000000";
--			ram(156) <= "00000000";
--			ram(157) <= "00000000";
--			ram(158) <= "00000000";
--			ram(159) <= "00000000";
--			ram(160) <= "00000000";
--			ram(161) <= "00000000";
--			ram(162) <= "00000000";
--			ram(163) <= "00000000";
--			ram(164) <= "00000000";
--			ram(165) <= "00000000";
--			ram(166) <= "00000000";
--			ram(167) <= "00000000";
--			ram(168) <= "00000000";
--			ram(169) <= "00000000";
--			ram(170) <= "00000000";
--			ram(171) <= "00000000";
--			ram(172) <= "00000000";
--			ram(173) <= "00000000";
--			ram(174) <= "00000000";
--			ram(175) <= "00000000";
--			ram(176) <= "00000000";
--			ram(177) <= "00000000";
--			ram(178) <= "00000000";
--			ram(179) <= "00000000";
--			ram(180) <= "00000000";
--			ram(181) <= "00000000";
--			ram(182) <= "00000000";
--			ram(183) <= "00000000";
--			ram(184) <= "00000000";
--			ram(185) <= "00000000";
--			ram(186) <= "00000000";
--			ram(187) <= "00000000";
--			ram(188) <= "00000000";
--			ram(189) <= "00000000";
--			ram(190) <= "00000000";
--			ram(191) <= "00000000";
--			ram(192) <= "00000000";
--			ram(193) <= "00000000";
--			ram(194) <= "00000000";
--			ram(195) <= "00000000";
--			ram(196) <= "00000000";
--			ram(197) <= "00000000";
--			ram(198) <= "00000000";
--			ram(199) <= "00000000";
--			ram(200) <= "00000000";
--			ram(201) <= "00000000";
--			ram(202) <= "00000000";
--			ram(203) <= "00000000";
--			ram(204) <= "00000000";
--			ram(205) <= "00000000";
--			ram(206) <= "00000000";
--			ram(207) <= "00000000";
--			ram(208) <= "00000000";
--			ram(209) <= "00000000";
--			ram(210) <= "00000000";
--			ram(211) <= "00000000";
--			ram(212) <= "00000000";
--			ram(213) <= "00000000";
--			ram(214) <= "00000000";
--			ram(215) <= "00000000";
--			ram(216) <= "00000000";
--			ram(217) <= "00000000";
--			ram(218) <= "00000000";
--			ram(219) <= "00000000";
--			ram(220) <= "00000000";
--			ram(221) <= "00000000";
--			ram(222) <= "00000000";
--			ram(223) <= "00000000";
--			ram(224) <= "00000000";
--			ram(225) <= "00000000";
--			ram(226) <= "00000000";
--			ram(227) <= "00000000";
--			ram(228) <= "00000000";
--			ram(229) <= "00000000";
--			ram(230) <= "00000000";
--			ram(231) <= "00000000";
--			ram(232) <= "00000000";
--			ram(233) <= "00000000";
--			ram(234) <= "00000000";
--			ram(235) <= "00000000";
--			ram(236) <= "00000000";
--			ram(237) <= "00000000";
--			ram(238) <= "00000000";
--			ram(239) <= "00000000";
--			ram(240) <= "00000000";
--			ram(241) <= "00000000";
--			ram(242) <= "00000000";
--			ram(243) <= "00000000";
--			ram(244) <= "00000000";
--			ram(245) <= "00000000";
--			ram(246) <= "00000000";
--			ram(247) <= "00000000";
--			ram(248) <= "00000000";
--			ram(249) <= "00000000";
--			ram(250) <= "00000000";
--			ram(251) <= "00000000";
--			ram(252) <= "00000000";
--			ram(253) <= "00000000";
--			ram(254) <= "00000000";
--			ram(255) <= "00000000";
--			ram(256) <= "00000000";
--			ram(257) <= "00000000";
--			ram(258) <= "00000000";
--			ram(259) <= "00000000";
--			ram(260) <= "00000000";
--			ram(261) <= "00000000";
--			ram(262) <= "00000000";
--			ram(263) <= "00000000";
--			ram(264) <= "00000000";
--			ram(265) <= "00000000";
--			ram(266) <= "00000000";
--			ram(267) <= "00000000";
--			ram(268) <= "00000000";
--			ram(269) <= "00000000";
--			ram(270) <= "00000000";
--			ram(271) <= "00000000";
--			ram(272) <= "00000000";
--			ram(273) <= "00000000";
--			ram(274) <= "00000000";
--			ram(275) <= "00000000";
--			ram(276) <= "00000000";
--			ram(277) <= "00000000";
--			ram(278) <= "00000000";
--			ram(279) <= "00000000";
--			ram(280) <= "00000000";
--			ram(281) <= "00000000";
--			ram(282) <= "00000000";
--			ram(283) <= "00000000";
--			ram(284) <= "00000000";
--			ram(285) <= "00000000";
--			ram(286) <= "00000000";
--			ram(287) <= "00000000";
--			ram(288) <= "00000000";
--			ram(289) <= "00000000";
--			ram(290) <= "00000000";
--			ram(291) <= "00000000";
--			ram(292) <= "00000000";
--			ram(293) <= "00000000";
--			ram(294) <= "00000000";
--			ram(295) <= "00000000";
--			ram(296) <= "00000000";
--			ram(297) <= "00000000";
--			ram(298) <= "00000000";
--			ram(299) <= "00000000";
--			ram(300) <= "00000000";
--			ram(301) <= "00000000";
--			ram(302) <= "00000000";
--			ram(303) <= "00000000";
--			ram(304) <= "00000000";
--			ram(305) <= "00000000";
--			ram(306) <= "00000000";
--			ram(307) <= "00000000";
--			ram(308) <= "00000000";
--			ram(309) <= "00000000";
--			ram(310) <= "00000000";
--			ram(311) <= "00000000";
--			ram(312) <= "00000000";
--			ram(313) <= "00000000";
--			ram(314) <= "00000000";
--			ram(315) <= "00000000";
--			ram(316) <= "00000000";
--			ram(317) <= "00000000";
--			ram(318) <= "00000000";
--			ram(319) <= "00000000";
--			ram(320) <= "00000000";
--			ram(321) <= "00000000";
--			ram(322) <= "00000000";
--			ram(323) <= "00000000";
--			ram(324) <= "00000000";
--			ram(325) <= "00000000";
--			ram(326) <= "00000000";
--			ram(327) <= "00000000";
--			ram(328) <= "00000000";
--			ram(329) <= "00000000";
--			ram(330) <= "00000000";
--			ram(331) <= "00000000";
--			ram(332) <= "00000000";
--			ram(333) <= "00000000";
--			ram(334) <= "00000000";
--			ram(335) <= "00000000";
--			ram(336) <= "00000000";
--			ram(337) <= "00000000";
--			ram(338) <= "00000000";
--			ram(339) <= "00000000";
--			ram(340) <= "00000000";
--			ram(341) <= "00000000";
--			ram(342) <= "00000000";
--			ram(343) <= "00000000";
--			ram(344) <= "00000000";
--			ram(345) <= "00000000";
--			ram(346) <= "00000000";
--			ram(347) <= "00000000";
--			ram(348) <= "00000000";
--			ram(349) <= "00000000";
--			ram(350) <= "00000000";
--			ram(351) <= "00000000";
--			ram(352) <= "00000000";
--			ram(353) <= "00000000";
--			ram(354) <= "00000000";
--			ram(355) <= "00000000";
--			ram(356) <= "00000000";
--			ram(357) <= "00000000";
--			ram(358) <= "00000000";
--			ram(359) <= "00000000";
--			ram(360) <= "00000000";
--			ram(361) <= "00000000";
--			ram(362) <= "00000000";
--			ram(363) <= "00000000";
--			ram(364) <= "00000000";
--			ram(365) <= "00000000";
--			ram(366) <= "00000000";
--			ram(367) <= "00000000";
--			ram(368) <= "00000000";
--			ram(369) <= "00000000";
--			ram(370) <= "00000000";
--			ram(371) <= "00000000";
--			ram(372) <= "00000000";
--			ram(373) <= "00000000";
--			ram(374) <= "00000000";
--			ram(375) <= "00000000";
--			ram(376) <= "00000000";
--			ram(377) <= "00000000";
--			ram(378) <= "00000000";
--			ram(379) <= "00000000";
--			ram(380) <= "00000000";
--			ram(381) <= "00000000";
--			ram(382) <= "00000000";
--			ram(383) <= "00000000";
--			ram(384) <= "00000000";
--			ram(385) <= "00000000";
--			ram(386) <= "00000000";
--			ram(387) <= "00000000";
--			ram(388) <= "00000000";
--			ram(389) <= "00000000";
--			ram(390) <= "00000000";
--			ram(391) <= "00000000";
--			ram(392) <= "00000000";
--			ram(393) <= "00000000";
--			ram(394) <= "00000000";
--			ram(395) <= "00000000";
--			ram(396) <= "00000000";
--			ram(397) <= "00000000";
--			ram(398) <= "00000000";
--			ram(399) <= "00000000";
--			ram(400) <= "00000000";
--			ram(401) <= "00000000";
--			ram(402) <= "00000000";
--			ram(403) <= "00000000";
--			ram(404) <= "00000000";
--			ram(405) <= "00000000";
--			ram(406) <= "00000000";
--			ram(407) <= "00000000";
--			ram(408) <= "00000000";
--			ram(409) <= "00000000";
--			ram(410) <= "00000000";
--			ram(411) <= "00000000";
--			ram(412) <= "00000000";
--			ram(413) <= "00000000";
--			ram(414) <= "00000000";
--			ram(415) <= "00000000";
--			ram(416) <= "00000000";
--			ram(417) <= "00000000";
--			ram(418) <= "00000000";
--			ram(419) <= "00000000";
--			ram(420) <= "00000000";
--			ram(421) <= "00000000";
--			ram(422) <= "00000000";
--			ram(423) <= "00000000";
--			ram(424) <= "00000000";
--			ram(425) <= "00000000";
--			ram(426) <= "00000000";
--			ram(427) <= "00000000";
--			ram(428) <= "00000000";
--			ram(429) <= "00000000";
--			ram(430) <= "00000000";
--			ram(431) <= "00000000";
--			ram(432) <= "00000000";
--			ram(433) <= "00000000";
--			ram(434) <= "00000000";
--			ram(435) <= "00000000";
--			ram(436) <= "00000000";
--			ram(437) <= "00000000";
--			ram(438) <= "00000000";
--			ram(439) <= "00000000";
--			ram(440) <= "00000000";
--			ram(441) <= "00000000";
--			ram(442) <= "00000000";
--			ram(443) <= "00000000";
--			ram(444) <= "00000000";
--			ram(445) <= "00000000";
--			ram(446) <= "00000000";
--			ram(447) <= "00000000";
--			ram(448) <= "00000000";
--			ram(449) <= "00000000";
--			ram(450) <= "00000000";
--			ram(451) <= "00000000";
--			ram(452) <= "00000000";
--			ram(453) <= "00000000";
--			ram(454) <= "00000000";
--			ram(455) <= "00000000";
--			ram(456) <= "00000000";
--			ram(457) <= "00000000";
--			ram(458) <= "00000000";
--			ram(459) <= "00000000";
--			ram(460) <= "00000000";
--			ram(461) <= "00000000";
--			ram(462) <= "00000000";
--			ram(463) <= "00000000";
--			ram(464) <= "00000000";
--			ram(465) <= "00000000";
--			ram(466) <= "00000000";
--			ram(467) <= "00000000";
--			ram(468) <= "00000000";
--			ram(469) <= "00000000";
--			ram(470) <= "00000000";
--			ram(471) <= "00000000";
--			ram(472) <= "00000000";
--			ram(473) <= "00000000";
--			ram(474) <= "00000000";
--			ram(475) <= "00000000";
--			ram(476) <= "00000000";
--			ram(477) <= "00000000";
--			ram(478) <= "00000000";
--			ram(479) <= "00000000";
--			ram(480) <= "00000000";
--			ram(481) <= "00000000";
--			ram(482) <= "00000000";
--			ram(483) <= "00000000";
--			ram(484) <= "00000000";
--			ram(485) <= "00000000";
--			ram(486) <= "00000000";
--			ram(487) <= "00000000";
--			ram(488) <= "00000000";
--			ram(489) <= "00000000";
--			ram(490) <= "00000000";
--			ram(491) <= "00000000";
--			ram(492) <= "00000000";
--			ram(493) <= "00000000";
--			ram(494) <= "00000000";
--			ram(495) <= "00000000";
--			ram(496) <= "00000000";
--			ram(497) <= "00000000";
--			ram(498) <= "00000000";
--			ram(499) <= "00000000";
--			ram(500) <= "00000000";
--			ram(501) <= "00000000";
--			ram(502) <= "00000000";
--			ram(503) <= "00000000";
--			ram(504) <= "00000000";
--			ram(505) <= "00000000";
--			ram(506) <= "00000000";
--			ram(507) <= "00000000";
--			ram(508) <= "00000000";
--			ram(509) <= "00000000";
--			ram(510) <= "00000000";
--			ram(511) <= "00000000";
--			ram(512) <= "00000000";
--			ram(513) <= "00000000";
--			ram(514) <= "00000000";
--			ram(515) <= "00000000";
--			ram(516) <= "00000000";
--			ram(517) <= "00000000";
--			ram(518) <= "00000000";
--			ram(519) <= "00000000";
--			ram(520) <= "00000000";
--			ram(521) <= "00000000";
--			ram(522) <= "00000000";
--			ram(523) <= "00000000";
--			ram(524) <= "00000000";
--			ram(525) <= "00000000";
--			ram(526) <= "00000000";
--			ram(527) <= "00000000";
--			ram(528) <= "00000000";
--			ram(529) <= "00000000";
--			ram(530) <= "00000000";
--			ram(531) <= "00000000";
--			ram(532) <= "00000000";
--			ram(533) <= "00000000";
--			ram(534) <= "00000000";
--			ram(535) <= "00000000";
--			ram(536) <= "00000000";
--			ram(537) <= "00000000";
--			ram(538) <= "00000000";
--			ram(539) <= "00000000";
--			ram(540) <= "00000000";
--			ram(541) <= "00000000";
--			ram(542) <= "00000000";
--			ram(543) <= "00000000";
--			ram(544) <= "00000000";
--			ram(545) <= "00000000";
--			ram(546) <= "00000000";
--			ram(547) <= "00000000";
--			ram(548) <= "00000000";
--			ram(549) <= "00000000";
--			ram(550) <= "00000000";
--			ram(551) <= "00000000";
--			ram(552) <= "00000000";
--			ram(553) <= "00000000";
--			ram(554) <= "00000000";
--			ram(555) <= "00000000";
--			ram(556) <= "00000000";
--			ram(557) <= "00000000";
--			ram(558) <= "00000000";
--			ram(559) <= "00000000";
--			ram(560) <= "00000000";
--			ram(561) <= "00000000";
--			ram(562) <= "00000000";
--			ram(563) <= "00000000";
--			ram(564) <= "00000000";
--			ram(565) <= "00000000";
--			ram(566) <= "00000000";
--			ram(567) <= "00000000";
--			ram(568) <= "00000000";
--			ram(569) <= "00000000";
--			ram(570) <= "00000000";
--			ram(571) <= "00000000";
--			ram(572) <= "00000000";
--			ram(573) <= "00000000";
--			ram(574) <= "00000000";
--			ram(575) <= "00000000";
--			ram(576) <= "00000000";
--			ram(577) <= "00000000";
--			ram(578) <= "00000000";
--			ram(579) <= "00000000";
--			ram(580) <= "00000000";
--			ram(581) <= "00000000";
--			ram(582) <= "00000000";
--			ram(583) <= "00000000";
--			ram(584) <= "00000000";
--			ram(585) <= "00000000";
--			ram(586) <= "00000000";
--			ram(587) <= "00000000";
--			ram(588) <= "00000000";
--			ram(589) <= "00000000";
--			ram(590) <= "00000000";
--			ram(591) <= "00000000";
--			ram(592) <= "00000000";
--			ram(593) <= "00000000";
--			ram(594) <= "00000000";
--			ram(595) <= "00000000";
--			ram(596) <= "00000000";
--			ram(597) <= "00000000";
--			ram(598) <= "00000000";
--			ram(599) <= "00000000";
--			ram(600) <= "00000000";
--			ram(601) <= "00000000";
--			ram(602) <= "00000000";
--			ram(603) <= "00000000";
--			ram(604) <= "00000000";
--			ram(605) <= "00000000";
--			ram(606) <= "00000000";
--			ram(607) <= "00000000";
--			ram(608) <= "00000000";
--			ram(609) <= "00000000";
--			ram(610) <= "00000000";
--			ram(611) <= "00000000";
--			ram(612) <= "00000000";
--			ram(613) <= "00000000";
--			ram(614) <= "00000000";
--			ram(615) <= "00000000";
--			ram(616) <= "00000000";
--			ram(617) <= "00000000";
--			ram(618) <= "00000000";
--			ram(619) <= "00000000";
--			ram(620) <= "00000000";
--			ram(621) <= "00000000";
--			ram(622) <= "00000000";
--			ram(623) <= "00000000";
--			ram(624) <= "00000000";
--			ram(625) <= "00000000";
--			ram(626) <= "00000000";
--			ram(627) <= "00000000";
--			ram(628) <= "00000000";
--			ram(629) <= "00000000";
--			ram(630) <= "00000000";
--			ram(631) <= "00000000";
--			ram(632) <= "00000000";
--			ram(633) <= "00000000";
--			ram(634) <= "00000000";
--			ram(635) <= "00000000";
--			ram(636) <= "00000000";
--			ram(637) <= "00000000";
--			ram(638) <= "00000000";
--			ram(639) <= "00000000";
--			ram(640) <= "00000000";
--			ram(641) <= "00000000";
--			ram(642) <= "00000000";
--			ram(643) <= "00000000";
--			ram(644) <= "00000000";
--			ram(645) <= "00000000";
--			ram(646) <= "00000000";
--			ram(647) <= "00000000";
--			ram(648) <= "00000000";
--			ram(649) <= "00000000";
--			ram(650) <= "00000000";
--			ram(651) <= "00000000";
--			ram(652) <= "00000000";
--			ram(653) <= "00000000";
--			ram(654) <= "00000000";
--			ram(655) <= "00000000";
--			ram(656) <= "00000000";
--			ram(657) <= "00000000";
--			ram(658) <= "00000000";
--			ram(659) <= "00000000";
--			ram(660) <= "00000000";
--			ram(661) <= "00000000";
--			ram(662) <= "00000000";
--			ram(663) <= "00000000";
--			ram(664) <= "00000000";
--			ram(665) <= "00000000";
--			ram(666) <= "00000000";
--			ram(667) <= "00000000";
--			ram(668) <= "00000000";
--			ram(669) <= "00000000";
--			ram(670) <= "00000000";
--			ram(671) <= "00000000";
--			ram(672) <= "00000000";
--			ram(673) <= "00000000";
--			ram(674) <= "00000000";
--			ram(675) <= "00000000";
--			ram(676) <= "00000000";
--			ram(677) <= "00000000";
--			ram(678) <= "00000000";
--			ram(679) <= "00000000";
--			ram(680) <= "00000000";
--			ram(681) <= "00000000";
--			ram(682) <= "00000000";
--			ram(683) <= "00000000";
--			ram(684) <= "00000000";
--			ram(685) <= "00000000";
--			ram(686) <= "00000000";
--			ram(687) <= "00000000";
--			ram(688) <= "00000000";
--			ram(689) <= "00000000";
--			ram(690) <= "00000000";
--			ram(691) <= "00000000";
--			ram(692) <= "00000000";
--			ram(693) <= "00000000";
--			ram(694) <= "00000000";
--			ram(695) <= "00000000";
--			ram(696) <= "00000000";
--			ram(697) <= "00000000";
--			ram(698) <= "00000000";
--			ram(699) <= "00000000";
--			ram(700) <= "00000000";
--			ram(701) <= "00000000";
--			ram(702) <= "00000000";
--			ram(703) <= "00000000";
--			ram(704) <= "00000000";
--			ram(705) <= "00000000";
--			ram(706) <= "00000000";
--			ram(707) <= "00000000";
--			ram(708) <= "00000000";
--			ram(709) <= "00000000";
--			ram(710) <= "00000000";
--			ram(711) <= "00000000";
--			ram(712) <= "00000000";
--			ram(713) <= "00000000";
--			ram(714) <= "00000000";
--			ram(715) <= "00000000";
--			ram(716) <= "00000000";
--			ram(717) <= "00000000";
--			ram(718) <= "00000000";
--			ram(719) <= "00000000";
--			ram(720) <= "00000000";
--			ram(721) <= "00000000";
--			ram(722) <= "00000000";
--			ram(723) <= "00000000";
--			ram(724) <= "00000000";
--			ram(725) <= "00000000";
--			ram(726) <= "00000000";
--			ram(727) <= "00000000";
--			ram(728) <= "00000000";
--			ram(729) <= "00000000";
--			ram(730) <= "00000000";
--			ram(731) <= "00000000";
--			ram(732) <= "00000000";
--			ram(733) <= "00000000";
--			ram(734) <= "00000000";
--			ram(735) <= "00000000";
--			ram(736) <= "00000000";
--			ram(737) <= "00000000";
--			ram(738) <= "00000000";
--			ram(739) <= "00000000";
--			ram(740) <= "00000000";
--			ram(741) <= "00000000";
--			ram(742) <= "00000000";
--			ram(743) <= "00000000";
--			ram(744) <= "00000000";
--			ram(745) <= "00000000";
--			ram(746) <= "00000000";
--			ram(747) <= "00000000";
--			ram(748) <= "00000000";
--			ram(749) <= "00000000";
--			ram(750) <= "00000000";
--			ram(751) <= "00000000";
--			ram(752) <= "00000000";
--			ram(753) <= "00000000";
--			ram(754) <= "00000000";
--			ram(755) <= "00000000";
--			ram(756) <= "00000000";
--			ram(757) <= "00000000";
--			ram(758) <= "00000000";
--			ram(759) <= "00000000";
--			ram(760) <= "00000000";
--			ram(761) <= "00000000";
--			ram(762) <= "00000000";
--			ram(763) <= "00000000";
--			ram(764) <= "00000000";
--			ram(765) <= "00000000";
--			ram(766) <= "00000000";
--			ram(767) <= "00000000";
--			ram(768) <= "00000000";
--			ram(769) <= "00000000";
--			ram(770) <= "00000000";
--			ram(771) <= "00000000";
--			ram(772) <= "00000000";
--			ram(773) <= "00000000";
--			ram(774) <= "00000000";
--			ram(775) <= "00000000";
--			ram(776) <= "00000000";
--			ram(777) <= "00000000";
--			ram(778) <= "00000000";
--			ram(779) <= "00000000";
--			ram(780) <= "00000000";
--			ram(781) <= "00000000";
--			ram(782) <= "00000000";
--			ram(783) <= "00000000";
--			ram(784) <= "00000000";
--			ram(785) <= "00000000";
--			ram(786) <= "00000000";
--			ram(787) <= "00000000";
--			ram(788) <= "00000000";
--			ram(789) <= "00000000";
--			ram(790) <= "00000000";
--			ram(791) <= "00000000";
--			ram(792) <= "00000000";
--			ram(793) <= "00000000";
--			ram(794) <= "00000000";
--			ram(795) <= "00000000";
--			ram(796) <= "00000000";
--			ram(797) <= "00000000";
--			ram(798) <= "00000000";
--			ram(799) <= "00000000";
--			ram(800) <= "00000000";
--			ram(801) <= "00000000";
--			ram(802) <= "00000000";
--			ram(803) <= "00000000";
--			ram(804) <= "00000000";
--			ram(805) <= "00000000";
--			ram(806) <= "00000000";
--			ram(807) <= "00000000";
--			ram(808) <= "00000000";
--			ram(809) <= "00000000";
--			ram(810) <= "00000000";
--			ram(811) <= "00000000";
--			ram(812) <= "00000000";
--			ram(813) <= "00000000";
--			ram(814) <= "00000000";
--			ram(815) <= "00000000";
--			ram(816) <= "00000000";
--			ram(817) <= "00000000";
--			ram(818) <= "00000000";
--			ram(819) <= "00000000";
--			ram(820) <= "00000000";
--			ram(821) <= "00000000";
--			ram(822) <= "00000000";
--			ram(823) <= "00000000";
--			ram(824) <= "00000000";
--			ram(825) <= "00000000";
--			ram(826) <= "00000000";
--			ram(827) <= "00000000";
--			ram(828) <= "00000000";
--			ram(829) <= "00000000";
--			ram(830) <= "00000000";
--			ram(831) <= "00000000";
--			ram(832) <= "00000000";
--			ram(833) <= "00000000";
--			ram(834) <= "00000000";
--			ram(835) <= "00000000";
--			ram(836) <= "00000000";
--			ram(837) <= "00000000";
--			ram(838) <= "00000000";
--			ram(839) <= "00000000";
--			ram(840) <= "00000000";
--			ram(841) <= "00000000";
--			ram(842) <= "00000000";
--			ram(843) <= "00000000";
--			ram(844) <= "00000000";
--			ram(845) <= "00000000";
--			ram(846) <= "00000000";
--			ram(847) <= "00000000";
--			ram(848) <= "00000000";
--			ram(849) <= "00000000";
--			ram(850) <= "00000000";
--			ram(851) <= "00000000";
--			ram(852) <= "00000000";
--			ram(853) <= "00000000";
--			ram(854) <= "00000000";
--			ram(855) <= "00000000";
--			ram(856) <= "00000000";
--			ram(857) <= "00000000";
--			ram(858) <= "00000000";
--			ram(859) <= "00000000";
--			ram(860) <= "00000000";
--			ram(861) <= "00000000";
--			ram(862) <= "00000000";
--			ram(863) <= "00000000";
--			ram(864) <= "00000000";
--			ram(865) <= "00000000";
--			ram(866) <= "00000000";
--			ram(867) <= "00000000";
--			ram(868) <= "00000000";
--			ram(869) <= "00000000";
--			ram(870) <= "00000000";
--			ram(871) <= "00000000";
--			ram(872) <= "00000000";
--			ram(873) <= "00000000";
--			ram(874) <= "00000000";
--			ram(875) <= "00000000";
--			ram(876) <= "00000000";
--			ram(877) <= "00000000";
--			ram(878) <= "00000000";
--			ram(879) <= "00000000";
--			ram(880) <= "00000000";
--			ram(881) <= "00000000";
--			ram(882) <= "00000000";
--			ram(883) <= "00000000";
--			ram(884) <= "00000000";
--			ram(885) <= "00000000";
--			ram(886) <= "00000000";
--			ram(887) <= "00000000";
--			ram(888) <= "00000000";
--			ram(889) <= "00000000";
--			ram(890) <= "00000000";
--			ram(891) <= "00000000";
--			ram(892) <= "00000000";
--			ram(893) <= "00000000";
--			ram(894) <= "00000000";
--			ram(895) <= "00000000";
--			ram(896) <= "00000000";
--			ram(897) <= "00000000";
--			ram(898) <= "00000000";
--			ram(899) <= "00000000";
--			ram(900) <= "00000000";
--			ram(901) <= "00000000";
--			ram(902) <= "00000000";
--			ram(903) <= "00000000";
--			ram(904) <= "00000000";
--			ram(905) <= "00000000";
--			ram(906) <= "00000000";
--			ram(907) <= "00000000";
--			ram(908) <= "00000000";
--			ram(909) <= "00000000";
--			ram(910) <= "00000000";
--			ram(911) <= "00000000";
--			ram(912) <= "00000000";
--			ram(913) <= "00000000";
--			ram(914) <= "00000000";
--			ram(915) <= "00000000";
--			ram(916) <= "00000000";
--			ram(917) <= "00000000";
--			ram(918) <= "00000000";
--			ram(919) <= "00000000";
--			ram(920) <= "00000000";
--			ram(921) <= "00000000";
--			ram(922) <= "00000000";
--			ram(923) <= "00000000";
--			ram(924) <= "00000000";
--			ram(925) <= "00000000";
--			ram(926) <= "00000000";
--			ram(927) <= "00000000";
--			ram(928) <= "00000000";
--			ram(929) <= "00000000";
--			ram(930) <= "00000000";
--			ram(931) <= "00000000";
--			ram(932) <= "00000000";
--			ram(933) <= "00000000";
--			ram(934) <= "00000000";
--			ram(935) <= "00000000";
--			ram(936) <= "00000000";
--			ram(937) <= "00000000";
--			ram(938) <= "00000000";
--			ram(939) <= "00000000";
--			ram(940) <= "00000000";
--			ram(941) <= "00000000";
--			ram(942) <= "00000000";
--			ram(943) <= "00000000";
--			ram(944) <= "00000000";
--			ram(945) <= "00000000";
--			ram(946) <= "00000000";
--			ram(947) <= "00000000";
--			ram(948) <= "00000000";
--			ram(949) <= "00000000";
--			ram(950) <= "00000000";
--			ram(951) <= "00000000";
--			ram(952) <= "00000000";
--			ram(953) <= "00000000";
--			ram(954) <= "00000000";
--			ram(955) <= "00000000";
--			ram(956) <= "00000000";
--			ram(957) <= "00000000";
--			ram(958) <= "00000000";
--			ram(959) <= "00000000";
--			ram(960) <= "00000000";
--			ram(961) <= "00000000";
--			ram(962) <= "00000000";
--			ram(963) <= "00000000";
--			ram(964) <= "00000000";
--			ram(965) <= "00000000";
--			ram(966) <= "00000000";
--			ram(967) <= "00000000";
--			ram(968) <= "00000000";
--			ram(969) <= "00000000";
--			ram(970) <= "00000000";
--			ram(971) <= "00000000";
--			ram(972) <= "00000000";
--			ram(973) <= "00000000";
--			ram(974) <= "00000000";
--			ram(975) <= "00000000";
--			ram(976) <= "00000000";
--			ram(977) <= "00000000";
--			ram(978) <= "00000000";
--			ram(979) <= "00000000";
--			ram(980) <= "00000000";
--			ram(981) <= "00000000";
--			ram(982) <= "00000000";
--			ram(983) <= "00000000";
--			ram(984) <= "00000000";
--			ram(985) <= "00000000";
--			ram(986) <= "00000000";
--			ram(987) <= "00000000";
--			ram(988) <= "00000000";
--			ram(989) <= "00000000";
--			ram(990) <= "00000000";
--			ram(991) <= "00000000";
--			ram(992) <= "00000000";
--			ram(993) <= "00000000";
--			ram(994) <= "00000000";
--			ram(995) <= "00000000";
--			ram(996) <= "00000000";
--			ram(997) <= "00000000";
--			ram(998) <= "00000000";
--			ram(999) <= "00000000";
--			ram(1000) <= "00000000";
--			ram(1001) <= "00000000";
--			ram(1002) <= "00000000";
--			ram(1003) <= "00000000";
--			ram(1004) <= "00000000";
--			ram(1005) <= "00000000";
--			ram(1006) <= "00000000";
--			ram(1007) <= "00000000";
--			ram(1008) <= "00000000";
--			ram(1009) <= "00000000";
--			ram(1010) <= "00000000";
--			ram(1011) <= "00000000";
--			ram(1012) <= "00000000";
--			ram(1013) <= "00000000";
--			ram(1014) <= "00000000";
--			ram(1015) <= "00000000";
--			ram(1016) <= "00000000";
--			ram(1017) <= "00000000";
--			ram(1018) <= "00000000";
--			ram(1019) <= "00000000";
--			ram(1020) <= "00000000";
--			ram(1021) <= "00000000";
--			ram(1022) <= "00000000";
--			ram(1023) <= "00000000";
			
		if (falling_edge(clk)) then
			var_addr := conv_integer(addr);
			if wr_en = '1' then
				ram(var_addr) <= data_in;
			end if;
				data_out <= ram(var_addr);
		end if;			
	end process;
end Behavioral;

